magic
tech sky130A
magscale 1 2
timestamp 1655310764
<< obsli1 >>
rect 1104 2159 248860 247537
<< obsm1 >>
rect 198 2128 249674 247568
<< metal2 >>
rect 4434 249200 4490 250000
rect 13358 249200 13414 250000
rect 22282 249200 22338 250000
rect 31206 249200 31262 250000
rect 40130 249200 40186 250000
rect 49054 249200 49110 250000
rect 57978 249200 58034 250000
rect 66902 249200 66958 250000
rect 75826 249200 75882 250000
rect 84750 249200 84806 250000
rect 93674 249200 93730 250000
rect 102598 249200 102654 250000
rect 111522 249200 111578 250000
rect 120446 249200 120502 250000
rect 129370 249200 129426 250000
rect 138294 249200 138350 250000
rect 147218 249200 147274 250000
rect 156142 249200 156198 250000
rect 165066 249200 165122 250000
rect 173990 249200 174046 250000
rect 182914 249200 182970 250000
rect 191838 249200 191894 250000
rect 200762 249200 200818 250000
rect 209686 249200 209742 250000
rect 218610 249200 218666 250000
rect 227534 249200 227590 250000
rect 236458 249200 236514 250000
rect 245382 249200 245438 250000
rect 202 0 258 800
rect 662 0 718 800
rect 1214 0 1270 800
rect 1674 0 1730 800
rect 2226 0 2282 800
rect 2686 0 2742 800
rect 3238 0 3294 800
rect 3698 0 3754 800
rect 4250 0 4306 800
rect 4710 0 4766 800
rect 5262 0 5318 800
rect 5722 0 5778 800
rect 6274 0 6330 800
rect 6734 0 6790 800
rect 7286 0 7342 800
rect 7838 0 7894 800
rect 8298 0 8354 800
rect 8850 0 8906 800
rect 9310 0 9366 800
rect 9862 0 9918 800
rect 10322 0 10378 800
rect 10874 0 10930 800
rect 11334 0 11390 800
rect 11886 0 11942 800
rect 12346 0 12402 800
rect 12898 0 12954 800
rect 13358 0 13414 800
rect 13910 0 13966 800
rect 14370 0 14426 800
rect 14922 0 14978 800
rect 15474 0 15530 800
rect 15934 0 15990 800
rect 16486 0 16542 800
rect 16946 0 17002 800
rect 17498 0 17554 800
rect 17958 0 18014 800
rect 18510 0 18566 800
rect 18970 0 19026 800
rect 19522 0 19578 800
rect 19982 0 20038 800
rect 20534 0 20590 800
rect 20994 0 21050 800
rect 21546 0 21602 800
rect 22006 0 22062 800
rect 22558 0 22614 800
rect 23110 0 23166 800
rect 23570 0 23626 800
rect 24122 0 24178 800
rect 24582 0 24638 800
rect 25134 0 25190 800
rect 25594 0 25650 800
rect 26146 0 26202 800
rect 26606 0 26662 800
rect 27158 0 27214 800
rect 27618 0 27674 800
rect 28170 0 28226 800
rect 28630 0 28686 800
rect 29182 0 29238 800
rect 29642 0 29698 800
rect 30194 0 30250 800
rect 30746 0 30802 800
rect 31206 0 31262 800
rect 31758 0 31814 800
rect 32218 0 32274 800
rect 32770 0 32826 800
rect 33230 0 33286 800
rect 33782 0 33838 800
rect 34242 0 34298 800
rect 34794 0 34850 800
rect 35254 0 35310 800
rect 35806 0 35862 800
rect 36266 0 36322 800
rect 36818 0 36874 800
rect 37278 0 37334 800
rect 37830 0 37886 800
rect 38382 0 38438 800
rect 38842 0 38898 800
rect 39394 0 39450 800
rect 39854 0 39910 800
rect 40406 0 40462 800
rect 40866 0 40922 800
rect 41418 0 41474 800
rect 41878 0 41934 800
rect 42430 0 42486 800
rect 42890 0 42946 800
rect 43442 0 43498 800
rect 43902 0 43958 800
rect 44454 0 44510 800
rect 44914 0 44970 800
rect 45466 0 45522 800
rect 46018 0 46074 800
rect 46478 0 46534 800
rect 47030 0 47086 800
rect 47490 0 47546 800
rect 48042 0 48098 800
rect 48502 0 48558 800
rect 49054 0 49110 800
rect 49514 0 49570 800
rect 50066 0 50122 800
rect 50526 0 50582 800
rect 51078 0 51134 800
rect 51538 0 51594 800
rect 52090 0 52146 800
rect 52550 0 52606 800
rect 53102 0 53158 800
rect 53654 0 53710 800
rect 54114 0 54170 800
rect 54666 0 54722 800
rect 55126 0 55182 800
rect 55678 0 55734 800
rect 56138 0 56194 800
rect 56690 0 56746 800
rect 57150 0 57206 800
rect 57702 0 57758 800
rect 58162 0 58218 800
rect 58714 0 58770 800
rect 59174 0 59230 800
rect 59726 0 59782 800
rect 60186 0 60242 800
rect 60738 0 60794 800
rect 61290 0 61346 800
rect 61750 0 61806 800
rect 62302 0 62358 800
rect 62762 0 62818 800
rect 63314 0 63370 800
rect 63774 0 63830 800
rect 64326 0 64382 800
rect 64786 0 64842 800
rect 65338 0 65394 800
rect 65798 0 65854 800
rect 66350 0 66406 800
rect 66810 0 66866 800
rect 67362 0 67418 800
rect 67822 0 67878 800
rect 68374 0 68430 800
rect 68926 0 68982 800
rect 69386 0 69442 800
rect 69938 0 69994 800
rect 70398 0 70454 800
rect 70950 0 71006 800
rect 71410 0 71466 800
rect 71962 0 72018 800
rect 72422 0 72478 800
rect 72974 0 73030 800
rect 73434 0 73490 800
rect 73986 0 74042 800
rect 74446 0 74502 800
rect 74998 0 75054 800
rect 75458 0 75514 800
rect 76010 0 76066 800
rect 76562 0 76618 800
rect 77022 0 77078 800
rect 77574 0 77630 800
rect 78034 0 78090 800
rect 78586 0 78642 800
rect 79046 0 79102 800
rect 79598 0 79654 800
rect 80058 0 80114 800
rect 80610 0 80666 800
rect 81070 0 81126 800
rect 81622 0 81678 800
rect 82082 0 82138 800
rect 82634 0 82690 800
rect 83094 0 83150 800
rect 83646 0 83702 800
rect 84198 0 84254 800
rect 84658 0 84714 800
rect 85210 0 85266 800
rect 85670 0 85726 800
rect 86222 0 86278 800
rect 86682 0 86738 800
rect 87234 0 87290 800
rect 87694 0 87750 800
rect 88246 0 88302 800
rect 88706 0 88762 800
rect 89258 0 89314 800
rect 89718 0 89774 800
rect 90270 0 90326 800
rect 90730 0 90786 800
rect 91282 0 91338 800
rect 91834 0 91890 800
rect 92294 0 92350 800
rect 92846 0 92902 800
rect 93306 0 93362 800
rect 93858 0 93914 800
rect 94318 0 94374 800
rect 94870 0 94926 800
rect 95330 0 95386 800
rect 95882 0 95938 800
rect 96342 0 96398 800
rect 96894 0 96950 800
rect 97354 0 97410 800
rect 97906 0 97962 800
rect 98366 0 98422 800
rect 98918 0 98974 800
rect 99470 0 99526 800
rect 99930 0 99986 800
rect 100482 0 100538 800
rect 100942 0 100998 800
rect 101494 0 101550 800
rect 101954 0 102010 800
rect 102506 0 102562 800
rect 102966 0 103022 800
rect 103518 0 103574 800
rect 103978 0 104034 800
rect 104530 0 104586 800
rect 104990 0 105046 800
rect 105542 0 105598 800
rect 106002 0 106058 800
rect 106554 0 106610 800
rect 107106 0 107162 800
rect 107566 0 107622 800
rect 108118 0 108174 800
rect 108578 0 108634 800
rect 109130 0 109186 800
rect 109590 0 109646 800
rect 110142 0 110198 800
rect 110602 0 110658 800
rect 111154 0 111210 800
rect 111614 0 111670 800
rect 112166 0 112222 800
rect 112626 0 112682 800
rect 113178 0 113234 800
rect 113638 0 113694 800
rect 114190 0 114246 800
rect 114742 0 114798 800
rect 115202 0 115258 800
rect 115754 0 115810 800
rect 116214 0 116270 800
rect 116766 0 116822 800
rect 117226 0 117282 800
rect 117778 0 117834 800
rect 118238 0 118294 800
rect 118790 0 118846 800
rect 119250 0 119306 800
rect 119802 0 119858 800
rect 120262 0 120318 800
rect 120814 0 120870 800
rect 121274 0 121330 800
rect 121826 0 121882 800
rect 122378 0 122434 800
rect 122838 0 122894 800
rect 123390 0 123446 800
rect 123850 0 123906 800
rect 124402 0 124458 800
rect 124862 0 124918 800
rect 125414 0 125470 800
rect 125874 0 125930 800
rect 126426 0 126482 800
rect 126886 0 126942 800
rect 127438 0 127494 800
rect 127898 0 127954 800
rect 128450 0 128506 800
rect 129002 0 129058 800
rect 129462 0 129518 800
rect 130014 0 130070 800
rect 130474 0 130530 800
rect 131026 0 131082 800
rect 131486 0 131542 800
rect 132038 0 132094 800
rect 132498 0 132554 800
rect 133050 0 133106 800
rect 133510 0 133566 800
rect 134062 0 134118 800
rect 134522 0 134578 800
rect 135074 0 135130 800
rect 135534 0 135590 800
rect 136086 0 136142 800
rect 136638 0 136694 800
rect 137098 0 137154 800
rect 137650 0 137706 800
rect 138110 0 138166 800
rect 138662 0 138718 800
rect 139122 0 139178 800
rect 139674 0 139730 800
rect 140134 0 140190 800
rect 140686 0 140742 800
rect 141146 0 141202 800
rect 141698 0 141754 800
rect 142158 0 142214 800
rect 142710 0 142766 800
rect 143170 0 143226 800
rect 143722 0 143778 800
rect 144274 0 144330 800
rect 144734 0 144790 800
rect 145286 0 145342 800
rect 145746 0 145802 800
rect 146298 0 146354 800
rect 146758 0 146814 800
rect 147310 0 147366 800
rect 147770 0 147826 800
rect 148322 0 148378 800
rect 148782 0 148838 800
rect 149334 0 149390 800
rect 149794 0 149850 800
rect 150346 0 150402 800
rect 150806 0 150862 800
rect 151358 0 151414 800
rect 151910 0 151966 800
rect 152370 0 152426 800
rect 152922 0 152978 800
rect 153382 0 153438 800
rect 153934 0 153990 800
rect 154394 0 154450 800
rect 154946 0 155002 800
rect 155406 0 155462 800
rect 155958 0 156014 800
rect 156418 0 156474 800
rect 156970 0 157026 800
rect 157430 0 157486 800
rect 157982 0 158038 800
rect 158442 0 158498 800
rect 158994 0 159050 800
rect 159546 0 159602 800
rect 160006 0 160062 800
rect 160558 0 160614 800
rect 161018 0 161074 800
rect 161570 0 161626 800
rect 162030 0 162086 800
rect 162582 0 162638 800
rect 163042 0 163098 800
rect 163594 0 163650 800
rect 164054 0 164110 800
rect 164606 0 164662 800
rect 165066 0 165122 800
rect 165618 0 165674 800
rect 166078 0 166134 800
rect 166630 0 166686 800
rect 167182 0 167238 800
rect 167642 0 167698 800
rect 168194 0 168250 800
rect 168654 0 168710 800
rect 169206 0 169262 800
rect 169666 0 169722 800
rect 170218 0 170274 800
rect 170678 0 170734 800
rect 171230 0 171286 800
rect 171690 0 171746 800
rect 172242 0 172298 800
rect 172702 0 172758 800
rect 173254 0 173310 800
rect 173714 0 173770 800
rect 174266 0 174322 800
rect 174818 0 174874 800
rect 175278 0 175334 800
rect 175830 0 175886 800
rect 176290 0 176346 800
rect 176842 0 176898 800
rect 177302 0 177358 800
rect 177854 0 177910 800
rect 178314 0 178370 800
rect 178866 0 178922 800
rect 179326 0 179382 800
rect 179878 0 179934 800
rect 180338 0 180394 800
rect 180890 0 180946 800
rect 181350 0 181406 800
rect 181902 0 181958 800
rect 182454 0 182510 800
rect 182914 0 182970 800
rect 183466 0 183522 800
rect 183926 0 183982 800
rect 184478 0 184534 800
rect 184938 0 184994 800
rect 185490 0 185546 800
rect 185950 0 186006 800
rect 186502 0 186558 800
rect 186962 0 187018 800
rect 187514 0 187570 800
rect 187974 0 188030 800
rect 188526 0 188582 800
rect 188986 0 189042 800
rect 189538 0 189594 800
rect 190090 0 190146 800
rect 190550 0 190606 800
rect 191102 0 191158 800
rect 191562 0 191618 800
rect 192114 0 192170 800
rect 192574 0 192630 800
rect 193126 0 193182 800
rect 193586 0 193642 800
rect 194138 0 194194 800
rect 194598 0 194654 800
rect 195150 0 195206 800
rect 195610 0 195666 800
rect 196162 0 196218 800
rect 196622 0 196678 800
rect 197174 0 197230 800
rect 197726 0 197782 800
rect 198186 0 198242 800
rect 198738 0 198794 800
rect 199198 0 199254 800
rect 199750 0 199806 800
rect 200210 0 200266 800
rect 200762 0 200818 800
rect 201222 0 201278 800
rect 201774 0 201830 800
rect 202234 0 202290 800
rect 202786 0 202842 800
rect 203246 0 203302 800
rect 203798 0 203854 800
rect 204258 0 204314 800
rect 204810 0 204866 800
rect 205362 0 205418 800
rect 205822 0 205878 800
rect 206374 0 206430 800
rect 206834 0 206890 800
rect 207386 0 207442 800
rect 207846 0 207902 800
rect 208398 0 208454 800
rect 208858 0 208914 800
rect 209410 0 209466 800
rect 209870 0 209926 800
rect 210422 0 210478 800
rect 210882 0 210938 800
rect 211434 0 211490 800
rect 211894 0 211950 800
rect 212446 0 212502 800
rect 212998 0 213054 800
rect 213458 0 213514 800
rect 214010 0 214066 800
rect 214470 0 214526 800
rect 215022 0 215078 800
rect 215482 0 215538 800
rect 216034 0 216090 800
rect 216494 0 216550 800
rect 217046 0 217102 800
rect 217506 0 217562 800
rect 218058 0 218114 800
rect 218518 0 218574 800
rect 219070 0 219126 800
rect 219530 0 219586 800
rect 220082 0 220138 800
rect 220634 0 220690 800
rect 221094 0 221150 800
rect 221646 0 221702 800
rect 222106 0 222162 800
rect 222658 0 222714 800
rect 223118 0 223174 800
rect 223670 0 223726 800
rect 224130 0 224186 800
rect 224682 0 224738 800
rect 225142 0 225198 800
rect 225694 0 225750 800
rect 226154 0 226210 800
rect 226706 0 226762 800
rect 227166 0 227222 800
rect 227718 0 227774 800
rect 228270 0 228326 800
rect 228730 0 228786 800
rect 229282 0 229338 800
rect 229742 0 229798 800
rect 230294 0 230350 800
rect 230754 0 230810 800
rect 231306 0 231362 800
rect 231766 0 231822 800
rect 232318 0 232374 800
rect 232778 0 232834 800
rect 233330 0 233386 800
rect 233790 0 233846 800
rect 234342 0 234398 800
rect 234802 0 234858 800
rect 235354 0 235410 800
rect 235906 0 235962 800
rect 236366 0 236422 800
rect 236918 0 236974 800
rect 237378 0 237434 800
rect 237930 0 237986 800
rect 238390 0 238446 800
rect 238942 0 238998 800
rect 239402 0 239458 800
rect 239954 0 240010 800
rect 240414 0 240470 800
rect 240966 0 241022 800
rect 241426 0 241482 800
rect 241978 0 242034 800
rect 242438 0 242494 800
rect 242990 0 243046 800
rect 243542 0 243598 800
rect 244002 0 244058 800
rect 244554 0 244610 800
rect 245014 0 245070 800
rect 245566 0 245622 800
rect 246026 0 246082 800
rect 246578 0 246634 800
rect 247038 0 247094 800
rect 247590 0 247646 800
rect 248050 0 248106 800
rect 248602 0 248658 800
rect 249062 0 249118 800
rect 249614 0 249670 800
<< obsm2 >>
rect 204 249144 4378 249234
rect 4546 249144 13302 249234
rect 13470 249144 22226 249234
rect 22394 249144 31150 249234
rect 31318 249144 40074 249234
rect 40242 249144 48998 249234
rect 49166 249144 57922 249234
rect 58090 249144 66846 249234
rect 67014 249144 75770 249234
rect 75938 249144 84694 249234
rect 84862 249144 93618 249234
rect 93786 249144 102542 249234
rect 102710 249144 111466 249234
rect 111634 249144 120390 249234
rect 120558 249144 129314 249234
rect 129482 249144 138238 249234
rect 138406 249144 147162 249234
rect 147330 249144 156086 249234
rect 156254 249144 165010 249234
rect 165178 249144 173934 249234
rect 174102 249144 182858 249234
rect 183026 249144 191782 249234
rect 191950 249144 200706 249234
rect 200874 249144 209630 249234
rect 209798 249144 218554 249234
rect 218722 249144 227478 249234
rect 227646 249144 236402 249234
rect 236570 249144 245326 249234
rect 245494 249144 249668 249234
rect 204 856 249668 249144
rect 314 800 606 856
rect 774 800 1158 856
rect 1326 800 1618 856
rect 1786 800 2170 856
rect 2338 800 2630 856
rect 2798 800 3182 856
rect 3350 800 3642 856
rect 3810 800 4194 856
rect 4362 800 4654 856
rect 4822 800 5206 856
rect 5374 800 5666 856
rect 5834 800 6218 856
rect 6386 800 6678 856
rect 6846 800 7230 856
rect 7398 800 7782 856
rect 7950 800 8242 856
rect 8410 800 8794 856
rect 8962 800 9254 856
rect 9422 800 9806 856
rect 9974 800 10266 856
rect 10434 800 10818 856
rect 10986 800 11278 856
rect 11446 800 11830 856
rect 11998 800 12290 856
rect 12458 800 12842 856
rect 13010 800 13302 856
rect 13470 800 13854 856
rect 14022 800 14314 856
rect 14482 800 14866 856
rect 15034 800 15418 856
rect 15586 800 15878 856
rect 16046 800 16430 856
rect 16598 800 16890 856
rect 17058 800 17442 856
rect 17610 800 17902 856
rect 18070 800 18454 856
rect 18622 800 18914 856
rect 19082 800 19466 856
rect 19634 800 19926 856
rect 20094 800 20478 856
rect 20646 800 20938 856
rect 21106 800 21490 856
rect 21658 800 21950 856
rect 22118 800 22502 856
rect 22670 800 23054 856
rect 23222 800 23514 856
rect 23682 800 24066 856
rect 24234 800 24526 856
rect 24694 800 25078 856
rect 25246 800 25538 856
rect 25706 800 26090 856
rect 26258 800 26550 856
rect 26718 800 27102 856
rect 27270 800 27562 856
rect 27730 800 28114 856
rect 28282 800 28574 856
rect 28742 800 29126 856
rect 29294 800 29586 856
rect 29754 800 30138 856
rect 30306 800 30690 856
rect 30858 800 31150 856
rect 31318 800 31702 856
rect 31870 800 32162 856
rect 32330 800 32714 856
rect 32882 800 33174 856
rect 33342 800 33726 856
rect 33894 800 34186 856
rect 34354 800 34738 856
rect 34906 800 35198 856
rect 35366 800 35750 856
rect 35918 800 36210 856
rect 36378 800 36762 856
rect 36930 800 37222 856
rect 37390 800 37774 856
rect 37942 800 38326 856
rect 38494 800 38786 856
rect 38954 800 39338 856
rect 39506 800 39798 856
rect 39966 800 40350 856
rect 40518 800 40810 856
rect 40978 800 41362 856
rect 41530 800 41822 856
rect 41990 800 42374 856
rect 42542 800 42834 856
rect 43002 800 43386 856
rect 43554 800 43846 856
rect 44014 800 44398 856
rect 44566 800 44858 856
rect 45026 800 45410 856
rect 45578 800 45962 856
rect 46130 800 46422 856
rect 46590 800 46974 856
rect 47142 800 47434 856
rect 47602 800 47986 856
rect 48154 800 48446 856
rect 48614 800 48998 856
rect 49166 800 49458 856
rect 49626 800 50010 856
rect 50178 800 50470 856
rect 50638 800 51022 856
rect 51190 800 51482 856
rect 51650 800 52034 856
rect 52202 800 52494 856
rect 52662 800 53046 856
rect 53214 800 53598 856
rect 53766 800 54058 856
rect 54226 800 54610 856
rect 54778 800 55070 856
rect 55238 800 55622 856
rect 55790 800 56082 856
rect 56250 800 56634 856
rect 56802 800 57094 856
rect 57262 800 57646 856
rect 57814 800 58106 856
rect 58274 800 58658 856
rect 58826 800 59118 856
rect 59286 800 59670 856
rect 59838 800 60130 856
rect 60298 800 60682 856
rect 60850 800 61234 856
rect 61402 800 61694 856
rect 61862 800 62246 856
rect 62414 800 62706 856
rect 62874 800 63258 856
rect 63426 800 63718 856
rect 63886 800 64270 856
rect 64438 800 64730 856
rect 64898 800 65282 856
rect 65450 800 65742 856
rect 65910 800 66294 856
rect 66462 800 66754 856
rect 66922 800 67306 856
rect 67474 800 67766 856
rect 67934 800 68318 856
rect 68486 800 68870 856
rect 69038 800 69330 856
rect 69498 800 69882 856
rect 70050 800 70342 856
rect 70510 800 70894 856
rect 71062 800 71354 856
rect 71522 800 71906 856
rect 72074 800 72366 856
rect 72534 800 72918 856
rect 73086 800 73378 856
rect 73546 800 73930 856
rect 74098 800 74390 856
rect 74558 800 74942 856
rect 75110 800 75402 856
rect 75570 800 75954 856
rect 76122 800 76506 856
rect 76674 800 76966 856
rect 77134 800 77518 856
rect 77686 800 77978 856
rect 78146 800 78530 856
rect 78698 800 78990 856
rect 79158 800 79542 856
rect 79710 800 80002 856
rect 80170 800 80554 856
rect 80722 800 81014 856
rect 81182 800 81566 856
rect 81734 800 82026 856
rect 82194 800 82578 856
rect 82746 800 83038 856
rect 83206 800 83590 856
rect 83758 800 84142 856
rect 84310 800 84602 856
rect 84770 800 85154 856
rect 85322 800 85614 856
rect 85782 800 86166 856
rect 86334 800 86626 856
rect 86794 800 87178 856
rect 87346 800 87638 856
rect 87806 800 88190 856
rect 88358 800 88650 856
rect 88818 800 89202 856
rect 89370 800 89662 856
rect 89830 800 90214 856
rect 90382 800 90674 856
rect 90842 800 91226 856
rect 91394 800 91778 856
rect 91946 800 92238 856
rect 92406 800 92790 856
rect 92958 800 93250 856
rect 93418 800 93802 856
rect 93970 800 94262 856
rect 94430 800 94814 856
rect 94982 800 95274 856
rect 95442 800 95826 856
rect 95994 800 96286 856
rect 96454 800 96838 856
rect 97006 800 97298 856
rect 97466 800 97850 856
rect 98018 800 98310 856
rect 98478 800 98862 856
rect 99030 800 99414 856
rect 99582 800 99874 856
rect 100042 800 100426 856
rect 100594 800 100886 856
rect 101054 800 101438 856
rect 101606 800 101898 856
rect 102066 800 102450 856
rect 102618 800 102910 856
rect 103078 800 103462 856
rect 103630 800 103922 856
rect 104090 800 104474 856
rect 104642 800 104934 856
rect 105102 800 105486 856
rect 105654 800 105946 856
rect 106114 800 106498 856
rect 106666 800 107050 856
rect 107218 800 107510 856
rect 107678 800 108062 856
rect 108230 800 108522 856
rect 108690 800 109074 856
rect 109242 800 109534 856
rect 109702 800 110086 856
rect 110254 800 110546 856
rect 110714 800 111098 856
rect 111266 800 111558 856
rect 111726 800 112110 856
rect 112278 800 112570 856
rect 112738 800 113122 856
rect 113290 800 113582 856
rect 113750 800 114134 856
rect 114302 800 114686 856
rect 114854 800 115146 856
rect 115314 800 115698 856
rect 115866 800 116158 856
rect 116326 800 116710 856
rect 116878 800 117170 856
rect 117338 800 117722 856
rect 117890 800 118182 856
rect 118350 800 118734 856
rect 118902 800 119194 856
rect 119362 800 119746 856
rect 119914 800 120206 856
rect 120374 800 120758 856
rect 120926 800 121218 856
rect 121386 800 121770 856
rect 121938 800 122322 856
rect 122490 800 122782 856
rect 122950 800 123334 856
rect 123502 800 123794 856
rect 123962 800 124346 856
rect 124514 800 124806 856
rect 124974 800 125358 856
rect 125526 800 125818 856
rect 125986 800 126370 856
rect 126538 800 126830 856
rect 126998 800 127382 856
rect 127550 800 127842 856
rect 128010 800 128394 856
rect 128562 800 128946 856
rect 129114 800 129406 856
rect 129574 800 129958 856
rect 130126 800 130418 856
rect 130586 800 130970 856
rect 131138 800 131430 856
rect 131598 800 131982 856
rect 132150 800 132442 856
rect 132610 800 132994 856
rect 133162 800 133454 856
rect 133622 800 134006 856
rect 134174 800 134466 856
rect 134634 800 135018 856
rect 135186 800 135478 856
rect 135646 800 136030 856
rect 136198 800 136582 856
rect 136750 800 137042 856
rect 137210 800 137594 856
rect 137762 800 138054 856
rect 138222 800 138606 856
rect 138774 800 139066 856
rect 139234 800 139618 856
rect 139786 800 140078 856
rect 140246 800 140630 856
rect 140798 800 141090 856
rect 141258 800 141642 856
rect 141810 800 142102 856
rect 142270 800 142654 856
rect 142822 800 143114 856
rect 143282 800 143666 856
rect 143834 800 144218 856
rect 144386 800 144678 856
rect 144846 800 145230 856
rect 145398 800 145690 856
rect 145858 800 146242 856
rect 146410 800 146702 856
rect 146870 800 147254 856
rect 147422 800 147714 856
rect 147882 800 148266 856
rect 148434 800 148726 856
rect 148894 800 149278 856
rect 149446 800 149738 856
rect 149906 800 150290 856
rect 150458 800 150750 856
rect 150918 800 151302 856
rect 151470 800 151854 856
rect 152022 800 152314 856
rect 152482 800 152866 856
rect 153034 800 153326 856
rect 153494 800 153878 856
rect 154046 800 154338 856
rect 154506 800 154890 856
rect 155058 800 155350 856
rect 155518 800 155902 856
rect 156070 800 156362 856
rect 156530 800 156914 856
rect 157082 800 157374 856
rect 157542 800 157926 856
rect 158094 800 158386 856
rect 158554 800 158938 856
rect 159106 800 159490 856
rect 159658 800 159950 856
rect 160118 800 160502 856
rect 160670 800 160962 856
rect 161130 800 161514 856
rect 161682 800 161974 856
rect 162142 800 162526 856
rect 162694 800 162986 856
rect 163154 800 163538 856
rect 163706 800 163998 856
rect 164166 800 164550 856
rect 164718 800 165010 856
rect 165178 800 165562 856
rect 165730 800 166022 856
rect 166190 800 166574 856
rect 166742 800 167126 856
rect 167294 800 167586 856
rect 167754 800 168138 856
rect 168306 800 168598 856
rect 168766 800 169150 856
rect 169318 800 169610 856
rect 169778 800 170162 856
rect 170330 800 170622 856
rect 170790 800 171174 856
rect 171342 800 171634 856
rect 171802 800 172186 856
rect 172354 800 172646 856
rect 172814 800 173198 856
rect 173366 800 173658 856
rect 173826 800 174210 856
rect 174378 800 174762 856
rect 174930 800 175222 856
rect 175390 800 175774 856
rect 175942 800 176234 856
rect 176402 800 176786 856
rect 176954 800 177246 856
rect 177414 800 177798 856
rect 177966 800 178258 856
rect 178426 800 178810 856
rect 178978 800 179270 856
rect 179438 800 179822 856
rect 179990 800 180282 856
rect 180450 800 180834 856
rect 181002 800 181294 856
rect 181462 800 181846 856
rect 182014 800 182398 856
rect 182566 800 182858 856
rect 183026 800 183410 856
rect 183578 800 183870 856
rect 184038 800 184422 856
rect 184590 800 184882 856
rect 185050 800 185434 856
rect 185602 800 185894 856
rect 186062 800 186446 856
rect 186614 800 186906 856
rect 187074 800 187458 856
rect 187626 800 187918 856
rect 188086 800 188470 856
rect 188638 800 188930 856
rect 189098 800 189482 856
rect 189650 800 190034 856
rect 190202 800 190494 856
rect 190662 800 191046 856
rect 191214 800 191506 856
rect 191674 800 192058 856
rect 192226 800 192518 856
rect 192686 800 193070 856
rect 193238 800 193530 856
rect 193698 800 194082 856
rect 194250 800 194542 856
rect 194710 800 195094 856
rect 195262 800 195554 856
rect 195722 800 196106 856
rect 196274 800 196566 856
rect 196734 800 197118 856
rect 197286 800 197670 856
rect 197838 800 198130 856
rect 198298 800 198682 856
rect 198850 800 199142 856
rect 199310 800 199694 856
rect 199862 800 200154 856
rect 200322 800 200706 856
rect 200874 800 201166 856
rect 201334 800 201718 856
rect 201886 800 202178 856
rect 202346 800 202730 856
rect 202898 800 203190 856
rect 203358 800 203742 856
rect 203910 800 204202 856
rect 204370 800 204754 856
rect 204922 800 205306 856
rect 205474 800 205766 856
rect 205934 800 206318 856
rect 206486 800 206778 856
rect 206946 800 207330 856
rect 207498 800 207790 856
rect 207958 800 208342 856
rect 208510 800 208802 856
rect 208970 800 209354 856
rect 209522 800 209814 856
rect 209982 800 210366 856
rect 210534 800 210826 856
rect 210994 800 211378 856
rect 211546 800 211838 856
rect 212006 800 212390 856
rect 212558 800 212942 856
rect 213110 800 213402 856
rect 213570 800 213954 856
rect 214122 800 214414 856
rect 214582 800 214966 856
rect 215134 800 215426 856
rect 215594 800 215978 856
rect 216146 800 216438 856
rect 216606 800 216990 856
rect 217158 800 217450 856
rect 217618 800 218002 856
rect 218170 800 218462 856
rect 218630 800 219014 856
rect 219182 800 219474 856
rect 219642 800 220026 856
rect 220194 800 220578 856
rect 220746 800 221038 856
rect 221206 800 221590 856
rect 221758 800 222050 856
rect 222218 800 222602 856
rect 222770 800 223062 856
rect 223230 800 223614 856
rect 223782 800 224074 856
rect 224242 800 224626 856
rect 224794 800 225086 856
rect 225254 800 225638 856
rect 225806 800 226098 856
rect 226266 800 226650 856
rect 226818 800 227110 856
rect 227278 800 227662 856
rect 227830 800 228214 856
rect 228382 800 228674 856
rect 228842 800 229226 856
rect 229394 800 229686 856
rect 229854 800 230238 856
rect 230406 800 230698 856
rect 230866 800 231250 856
rect 231418 800 231710 856
rect 231878 800 232262 856
rect 232430 800 232722 856
rect 232890 800 233274 856
rect 233442 800 233734 856
rect 233902 800 234286 856
rect 234454 800 234746 856
rect 234914 800 235298 856
rect 235466 800 235850 856
rect 236018 800 236310 856
rect 236478 800 236862 856
rect 237030 800 237322 856
rect 237490 800 237874 856
rect 238042 800 238334 856
rect 238502 800 238886 856
rect 239054 800 239346 856
rect 239514 800 239898 856
rect 240066 800 240358 856
rect 240526 800 240910 856
rect 241078 800 241370 856
rect 241538 800 241922 856
rect 242090 800 242382 856
rect 242550 800 242934 856
rect 243102 800 243486 856
rect 243654 800 243946 856
rect 244114 800 244498 856
rect 244666 800 244958 856
rect 245126 800 245510 856
rect 245678 800 245970 856
rect 246138 800 246522 856
rect 246690 800 246982 856
rect 247150 800 247534 856
rect 247702 800 247994 856
rect 248162 800 248546 856
rect 248714 800 249006 856
rect 249174 800 249558 856
<< metal3 >>
rect 249200 247120 250000 247240
rect 0 246848 800 246968
rect 249200 241680 250000 241800
rect 0 240864 800 240984
rect 249200 236240 250000 236360
rect 0 234880 800 235000
rect 249200 230800 250000 230920
rect 0 228896 800 229016
rect 249200 225360 250000 225480
rect 0 223048 800 223168
rect 249200 219920 250000 220040
rect 0 217064 800 217184
rect 249200 214480 250000 214600
rect 0 211080 800 211200
rect 249200 209040 250000 209160
rect 0 205096 800 205216
rect 249200 203600 250000 203720
rect 0 199248 800 199368
rect 249200 198160 250000 198280
rect 0 193264 800 193384
rect 249200 192720 250000 192840
rect 0 187280 800 187400
rect 249200 187280 250000 187400
rect 249200 181840 250000 181960
rect 0 181296 800 181416
rect 249200 176400 250000 176520
rect 0 175448 800 175568
rect 249200 170960 250000 171080
rect 0 169464 800 169584
rect 249200 165520 250000 165640
rect 0 163480 800 163600
rect 249200 160080 250000 160200
rect 0 157496 800 157616
rect 249200 154640 250000 154760
rect 0 151648 800 151768
rect 249200 149200 250000 149320
rect 0 145664 800 145784
rect 249200 143760 250000 143880
rect 0 139680 800 139800
rect 249200 138320 250000 138440
rect 0 133696 800 133816
rect 249200 132880 250000 133000
rect 0 127848 800 127968
rect 249200 127576 250000 127696
rect 249200 122136 250000 122256
rect 0 121864 800 121984
rect 249200 116696 250000 116816
rect 0 115880 800 116000
rect 249200 111256 250000 111376
rect 0 109896 800 110016
rect 249200 105816 250000 105936
rect 0 103912 800 104032
rect 249200 100376 250000 100496
rect 0 98064 800 98184
rect 249200 94936 250000 95056
rect 0 92080 800 92200
rect 249200 89496 250000 89616
rect 0 86096 800 86216
rect 249200 84056 250000 84176
rect 0 80112 800 80232
rect 249200 78616 250000 78736
rect 0 74264 800 74384
rect 249200 73176 250000 73296
rect 0 68280 800 68400
rect 249200 67736 250000 67856
rect 0 62296 800 62416
rect 249200 62296 250000 62416
rect 249200 56856 250000 56976
rect 0 56312 800 56432
rect 249200 51416 250000 51536
rect 0 50464 800 50584
rect 249200 45976 250000 46096
rect 0 44480 800 44600
rect 249200 40536 250000 40656
rect 0 38496 800 38616
rect 249200 35096 250000 35216
rect 0 32512 800 32632
rect 249200 29656 250000 29776
rect 0 26664 800 26784
rect 249200 24216 250000 24336
rect 0 20680 800 20800
rect 249200 18776 250000 18896
rect 0 14696 800 14816
rect 249200 13336 250000 13456
rect 0 8712 800 8832
rect 249200 7896 250000 8016
rect 0 2864 800 2984
rect 249200 2592 250000 2712
<< obsm3 >>
rect 800 247320 249200 247553
rect 800 247048 249120 247320
rect 880 247040 249120 247048
rect 880 246768 249200 247040
rect 800 241880 249200 246768
rect 800 241600 249120 241880
rect 800 241064 249200 241600
rect 880 240784 249200 241064
rect 800 236440 249200 240784
rect 800 236160 249120 236440
rect 800 235080 249200 236160
rect 880 234800 249200 235080
rect 800 231000 249200 234800
rect 800 230720 249120 231000
rect 800 229096 249200 230720
rect 880 228816 249200 229096
rect 800 225560 249200 228816
rect 800 225280 249120 225560
rect 800 223248 249200 225280
rect 880 222968 249200 223248
rect 800 220120 249200 222968
rect 800 219840 249120 220120
rect 800 217264 249200 219840
rect 880 216984 249200 217264
rect 800 214680 249200 216984
rect 800 214400 249120 214680
rect 800 211280 249200 214400
rect 880 211000 249200 211280
rect 800 209240 249200 211000
rect 800 208960 249120 209240
rect 800 205296 249200 208960
rect 880 205016 249200 205296
rect 800 203800 249200 205016
rect 800 203520 249120 203800
rect 800 199448 249200 203520
rect 880 199168 249200 199448
rect 800 198360 249200 199168
rect 800 198080 249120 198360
rect 800 193464 249200 198080
rect 880 193184 249200 193464
rect 800 192920 249200 193184
rect 800 192640 249120 192920
rect 800 187480 249200 192640
rect 880 187200 249120 187480
rect 800 182040 249200 187200
rect 800 181760 249120 182040
rect 800 181496 249200 181760
rect 880 181216 249200 181496
rect 800 176600 249200 181216
rect 800 176320 249120 176600
rect 800 175648 249200 176320
rect 880 175368 249200 175648
rect 800 171160 249200 175368
rect 800 170880 249120 171160
rect 800 169664 249200 170880
rect 880 169384 249200 169664
rect 800 165720 249200 169384
rect 800 165440 249120 165720
rect 800 163680 249200 165440
rect 880 163400 249200 163680
rect 800 160280 249200 163400
rect 800 160000 249120 160280
rect 800 157696 249200 160000
rect 880 157416 249200 157696
rect 800 154840 249200 157416
rect 800 154560 249120 154840
rect 800 151848 249200 154560
rect 880 151568 249200 151848
rect 800 149400 249200 151568
rect 800 149120 249120 149400
rect 800 145864 249200 149120
rect 880 145584 249200 145864
rect 800 143960 249200 145584
rect 800 143680 249120 143960
rect 800 139880 249200 143680
rect 880 139600 249200 139880
rect 800 138520 249200 139600
rect 800 138240 249120 138520
rect 800 133896 249200 138240
rect 880 133616 249200 133896
rect 800 133080 249200 133616
rect 800 132800 249120 133080
rect 800 128048 249200 132800
rect 880 127776 249200 128048
rect 880 127768 249120 127776
rect 800 127496 249120 127768
rect 800 122336 249200 127496
rect 800 122064 249120 122336
rect 880 122056 249120 122064
rect 880 121784 249200 122056
rect 800 116896 249200 121784
rect 800 116616 249120 116896
rect 800 116080 249200 116616
rect 880 115800 249200 116080
rect 800 111456 249200 115800
rect 800 111176 249120 111456
rect 800 110096 249200 111176
rect 880 109816 249200 110096
rect 800 106016 249200 109816
rect 800 105736 249120 106016
rect 800 104112 249200 105736
rect 880 103832 249200 104112
rect 800 100576 249200 103832
rect 800 100296 249120 100576
rect 800 98264 249200 100296
rect 880 97984 249200 98264
rect 800 95136 249200 97984
rect 800 94856 249120 95136
rect 800 92280 249200 94856
rect 880 92000 249200 92280
rect 800 89696 249200 92000
rect 800 89416 249120 89696
rect 800 86296 249200 89416
rect 880 86016 249200 86296
rect 800 84256 249200 86016
rect 800 83976 249120 84256
rect 800 80312 249200 83976
rect 880 80032 249200 80312
rect 800 78816 249200 80032
rect 800 78536 249120 78816
rect 800 74464 249200 78536
rect 880 74184 249200 74464
rect 800 73376 249200 74184
rect 800 73096 249120 73376
rect 800 68480 249200 73096
rect 880 68200 249200 68480
rect 800 67936 249200 68200
rect 800 67656 249120 67936
rect 800 62496 249200 67656
rect 880 62216 249120 62496
rect 800 57056 249200 62216
rect 800 56776 249120 57056
rect 800 56512 249200 56776
rect 880 56232 249200 56512
rect 800 51616 249200 56232
rect 800 51336 249120 51616
rect 800 50664 249200 51336
rect 880 50384 249200 50664
rect 800 46176 249200 50384
rect 800 45896 249120 46176
rect 800 44680 249200 45896
rect 880 44400 249200 44680
rect 800 40736 249200 44400
rect 800 40456 249120 40736
rect 800 38696 249200 40456
rect 880 38416 249200 38696
rect 800 35296 249200 38416
rect 800 35016 249120 35296
rect 800 32712 249200 35016
rect 880 32432 249200 32712
rect 800 29856 249200 32432
rect 800 29576 249120 29856
rect 800 26864 249200 29576
rect 880 26584 249200 26864
rect 800 24416 249200 26584
rect 800 24136 249120 24416
rect 800 20880 249200 24136
rect 880 20600 249200 20880
rect 800 18976 249200 20600
rect 800 18696 249120 18976
rect 800 14896 249200 18696
rect 880 14616 249200 14896
rect 800 13536 249200 14616
rect 800 13256 249120 13536
rect 800 8912 249200 13256
rect 880 8632 249200 8912
rect 800 8096 249200 8632
rect 800 7816 249120 8096
rect 800 3064 249200 7816
rect 880 2792 249200 3064
rect 880 2784 249120 2792
rect 800 2512 249120 2784
rect 800 2143 249200 2512
<< metal4 >>
rect 4208 2128 4528 247568
rect 19568 2128 19888 247568
rect 34928 2128 35248 247568
rect 50288 2128 50608 247568
rect 65648 2128 65968 247568
rect 81008 2128 81328 247568
rect 96368 2128 96688 247568
rect 111728 2128 112048 247568
rect 127088 2128 127408 247568
rect 142448 2128 142768 247568
rect 157808 2128 158128 247568
rect 173168 2128 173488 247568
rect 188528 2128 188848 247568
rect 203888 2128 204208 247568
rect 219248 2128 219568 247568
rect 234608 2128 234928 247568
<< obsm4 >>
rect 87275 46683 96288 179757
rect 96768 46683 111648 179757
rect 112128 46683 127008 179757
rect 127488 46683 142368 179757
rect 142848 46683 157728 179757
rect 158208 46683 173088 179757
rect 173568 46683 188448 179757
rect 188928 46683 203808 179757
rect 204288 46683 219168 179757
rect 219648 46683 234528 179757
rect 235008 46683 238037 179757
<< labels >>
rlabel metal3 s 249200 2592 250000 2712 6 io_in[0]
port 1 nsew signal input
rlabel metal3 s 249200 165520 250000 165640 6 io_in[10]
port 2 nsew signal input
rlabel metal3 s 249200 181840 250000 181960 6 io_in[11]
port 3 nsew signal input
rlabel metal3 s 249200 198160 250000 198280 6 io_in[12]
port 4 nsew signal input
rlabel metal3 s 249200 214480 250000 214600 6 io_in[13]
port 5 nsew signal input
rlabel metal3 s 249200 230800 250000 230920 6 io_in[14]
port 6 nsew signal input
rlabel metal2 s 245382 249200 245438 250000 6 io_in[15]
port 7 nsew signal input
rlabel metal2 s 218610 249200 218666 250000 6 io_in[16]
port 8 nsew signal input
rlabel metal2 s 191838 249200 191894 250000 6 io_in[17]
port 9 nsew signal input
rlabel metal2 s 165066 249200 165122 250000 6 io_in[18]
port 10 nsew signal input
rlabel metal2 s 138294 249200 138350 250000 6 io_in[19]
port 11 nsew signal input
rlabel metal3 s 249200 18776 250000 18896 6 io_in[1]
port 12 nsew signal input
rlabel metal2 s 111522 249200 111578 250000 6 io_in[20]
port 13 nsew signal input
rlabel metal2 s 84750 249200 84806 250000 6 io_in[21]
port 14 nsew signal input
rlabel metal2 s 57978 249200 58034 250000 6 io_in[22]
port 15 nsew signal input
rlabel metal2 s 31206 249200 31262 250000 6 io_in[23]
port 16 nsew signal input
rlabel metal3 s 0 246848 800 246968 6 io_in[24]
port 17 nsew signal input
rlabel metal3 s 0 228896 800 229016 6 io_in[25]
port 18 nsew signal input
rlabel metal3 s 0 211080 800 211200 6 io_in[26]
port 19 nsew signal input
rlabel metal3 s 0 193264 800 193384 6 io_in[27]
port 20 nsew signal input
rlabel metal3 s 0 175448 800 175568 6 io_in[28]
port 21 nsew signal input
rlabel metal3 s 0 157496 800 157616 6 io_in[29]
port 22 nsew signal input
rlabel metal3 s 249200 35096 250000 35216 6 io_in[2]
port 23 nsew signal input
rlabel metal3 s 0 139680 800 139800 6 io_in[30]
port 24 nsew signal input
rlabel metal3 s 0 121864 800 121984 6 io_in[31]
port 25 nsew signal input
rlabel metal3 s 0 103912 800 104032 6 io_in[32]
port 26 nsew signal input
rlabel metal3 s 0 86096 800 86216 6 io_in[33]
port 27 nsew signal input
rlabel metal3 s 0 68280 800 68400 6 io_in[34]
port 28 nsew signal input
rlabel metal3 s 0 50464 800 50584 6 io_in[35]
port 29 nsew signal input
rlabel metal3 s 0 32512 800 32632 6 io_in[36]
port 30 nsew signal input
rlabel metal3 s 0 14696 800 14816 6 io_in[37]
port 31 nsew signal input
rlabel metal3 s 249200 51416 250000 51536 6 io_in[3]
port 32 nsew signal input
rlabel metal3 s 249200 67736 250000 67856 6 io_in[4]
port 33 nsew signal input
rlabel metal3 s 249200 84056 250000 84176 6 io_in[5]
port 34 nsew signal input
rlabel metal3 s 249200 100376 250000 100496 6 io_in[6]
port 35 nsew signal input
rlabel metal3 s 249200 116696 250000 116816 6 io_in[7]
port 36 nsew signal input
rlabel metal3 s 249200 132880 250000 133000 6 io_in[8]
port 37 nsew signal input
rlabel metal3 s 249200 149200 250000 149320 6 io_in[9]
port 38 nsew signal input
rlabel metal3 s 249200 13336 250000 13456 6 io_oeb[0]
port 39 nsew signal output
rlabel metal3 s 249200 176400 250000 176520 6 io_oeb[10]
port 40 nsew signal output
rlabel metal3 s 249200 192720 250000 192840 6 io_oeb[11]
port 41 nsew signal output
rlabel metal3 s 249200 209040 250000 209160 6 io_oeb[12]
port 42 nsew signal output
rlabel metal3 s 249200 225360 250000 225480 6 io_oeb[13]
port 43 nsew signal output
rlabel metal3 s 249200 241680 250000 241800 6 io_oeb[14]
port 44 nsew signal output
rlabel metal2 s 227534 249200 227590 250000 6 io_oeb[15]
port 45 nsew signal output
rlabel metal2 s 200762 249200 200818 250000 6 io_oeb[16]
port 46 nsew signal output
rlabel metal2 s 173990 249200 174046 250000 6 io_oeb[17]
port 47 nsew signal output
rlabel metal2 s 147218 249200 147274 250000 6 io_oeb[18]
port 48 nsew signal output
rlabel metal2 s 120446 249200 120502 250000 6 io_oeb[19]
port 49 nsew signal output
rlabel metal3 s 249200 29656 250000 29776 6 io_oeb[1]
port 50 nsew signal output
rlabel metal2 s 93674 249200 93730 250000 6 io_oeb[20]
port 51 nsew signal output
rlabel metal2 s 66902 249200 66958 250000 6 io_oeb[21]
port 52 nsew signal output
rlabel metal2 s 40130 249200 40186 250000 6 io_oeb[22]
port 53 nsew signal output
rlabel metal2 s 13358 249200 13414 250000 6 io_oeb[23]
port 54 nsew signal output
rlabel metal3 s 0 234880 800 235000 6 io_oeb[24]
port 55 nsew signal output
rlabel metal3 s 0 217064 800 217184 6 io_oeb[25]
port 56 nsew signal output
rlabel metal3 s 0 199248 800 199368 6 io_oeb[26]
port 57 nsew signal output
rlabel metal3 s 0 181296 800 181416 6 io_oeb[27]
port 58 nsew signal output
rlabel metal3 s 0 163480 800 163600 6 io_oeb[28]
port 59 nsew signal output
rlabel metal3 s 0 145664 800 145784 6 io_oeb[29]
port 60 nsew signal output
rlabel metal3 s 249200 45976 250000 46096 6 io_oeb[2]
port 61 nsew signal output
rlabel metal3 s 0 127848 800 127968 6 io_oeb[30]
port 62 nsew signal output
rlabel metal3 s 0 109896 800 110016 6 io_oeb[31]
port 63 nsew signal output
rlabel metal3 s 0 92080 800 92200 6 io_oeb[32]
port 64 nsew signal output
rlabel metal3 s 0 74264 800 74384 6 io_oeb[33]
port 65 nsew signal output
rlabel metal3 s 0 56312 800 56432 6 io_oeb[34]
port 66 nsew signal output
rlabel metal3 s 0 38496 800 38616 6 io_oeb[35]
port 67 nsew signal output
rlabel metal3 s 0 20680 800 20800 6 io_oeb[36]
port 68 nsew signal output
rlabel metal3 s 0 2864 800 2984 6 io_oeb[37]
port 69 nsew signal output
rlabel metal3 s 249200 62296 250000 62416 6 io_oeb[3]
port 70 nsew signal output
rlabel metal3 s 249200 78616 250000 78736 6 io_oeb[4]
port 71 nsew signal output
rlabel metal3 s 249200 94936 250000 95056 6 io_oeb[5]
port 72 nsew signal output
rlabel metal3 s 249200 111256 250000 111376 6 io_oeb[6]
port 73 nsew signal output
rlabel metal3 s 249200 127576 250000 127696 6 io_oeb[7]
port 74 nsew signal output
rlabel metal3 s 249200 143760 250000 143880 6 io_oeb[8]
port 75 nsew signal output
rlabel metal3 s 249200 160080 250000 160200 6 io_oeb[9]
port 76 nsew signal output
rlabel metal3 s 249200 7896 250000 8016 6 io_out[0]
port 77 nsew signal output
rlabel metal3 s 249200 170960 250000 171080 6 io_out[10]
port 78 nsew signal output
rlabel metal3 s 249200 187280 250000 187400 6 io_out[11]
port 79 nsew signal output
rlabel metal3 s 249200 203600 250000 203720 6 io_out[12]
port 80 nsew signal output
rlabel metal3 s 249200 219920 250000 220040 6 io_out[13]
port 81 nsew signal output
rlabel metal3 s 249200 236240 250000 236360 6 io_out[14]
port 82 nsew signal output
rlabel metal2 s 236458 249200 236514 250000 6 io_out[15]
port 83 nsew signal output
rlabel metal2 s 209686 249200 209742 250000 6 io_out[16]
port 84 nsew signal output
rlabel metal2 s 182914 249200 182970 250000 6 io_out[17]
port 85 nsew signal output
rlabel metal2 s 156142 249200 156198 250000 6 io_out[18]
port 86 nsew signal output
rlabel metal2 s 129370 249200 129426 250000 6 io_out[19]
port 87 nsew signal output
rlabel metal3 s 249200 24216 250000 24336 6 io_out[1]
port 88 nsew signal output
rlabel metal2 s 102598 249200 102654 250000 6 io_out[20]
port 89 nsew signal output
rlabel metal2 s 75826 249200 75882 250000 6 io_out[21]
port 90 nsew signal output
rlabel metal2 s 49054 249200 49110 250000 6 io_out[22]
port 91 nsew signal output
rlabel metal2 s 22282 249200 22338 250000 6 io_out[23]
port 92 nsew signal output
rlabel metal3 s 0 240864 800 240984 6 io_out[24]
port 93 nsew signal output
rlabel metal3 s 0 223048 800 223168 6 io_out[25]
port 94 nsew signal output
rlabel metal3 s 0 205096 800 205216 6 io_out[26]
port 95 nsew signal output
rlabel metal3 s 0 187280 800 187400 6 io_out[27]
port 96 nsew signal output
rlabel metal3 s 0 169464 800 169584 6 io_out[28]
port 97 nsew signal output
rlabel metal3 s 0 151648 800 151768 6 io_out[29]
port 98 nsew signal output
rlabel metal3 s 249200 40536 250000 40656 6 io_out[2]
port 99 nsew signal output
rlabel metal3 s 0 133696 800 133816 6 io_out[30]
port 100 nsew signal output
rlabel metal3 s 0 115880 800 116000 6 io_out[31]
port 101 nsew signal output
rlabel metal3 s 0 98064 800 98184 6 io_out[32]
port 102 nsew signal output
rlabel metal3 s 0 80112 800 80232 6 io_out[33]
port 103 nsew signal output
rlabel metal3 s 0 62296 800 62416 6 io_out[34]
port 104 nsew signal output
rlabel metal3 s 0 44480 800 44600 6 io_out[35]
port 105 nsew signal output
rlabel metal3 s 0 26664 800 26784 6 io_out[36]
port 106 nsew signal output
rlabel metal3 s 0 8712 800 8832 6 io_out[37]
port 107 nsew signal output
rlabel metal3 s 249200 56856 250000 56976 6 io_out[3]
port 108 nsew signal output
rlabel metal3 s 249200 73176 250000 73296 6 io_out[4]
port 109 nsew signal output
rlabel metal3 s 249200 89496 250000 89616 6 io_out[5]
port 110 nsew signal output
rlabel metal3 s 249200 105816 250000 105936 6 io_out[6]
port 111 nsew signal output
rlabel metal3 s 249200 122136 250000 122256 6 io_out[7]
port 112 nsew signal output
rlabel metal3 s 249200 138320 250000 138440 6 io_out[8]
port 113 nsew signal output
rlabel metal3 s 249200 154640 250000 154760 6 io_out[9]
port 114 nsew signal output
rlabel metal2 s 249614 0 249670 800 6 irq[0]
port 115 nsew signal output
rlabel metal3 s 249200 247120 250000 247240 6 irq[1]
port 116 nsew signal output
rlabel metal2 s 4434 249200 4490 250000 6 irq[2]
port 117 nsew signal output
rlabel metal2 s 54114 0 54170 800 6 la_data_in[0]
port 118 nsew signal input
rlabel metal2 s 206834 0 206890 800 6 la_data_in[100]
port 119 nsew signal input
rlabel metal2 s 208398 0 208454 800 6 la_data_in[101]
port 120 nsew signal input
rlabel metal2 s 209870 0 209926 800 6 la_data_in[102]
port 121 nsew signal input
rlabel metal2 s 211434 0 211490 800 6 la_data_in[103]
port 122 nsew signal input
rlabel metal2 s 212998 0 213054 800 6 la_data_in[104]
port 123 nsew signal input
rlabel metal2 s 214470 0 214526 800 6 la_data_in[105]
port 124 nsew signal input
rlabel metal2 s 216034 0 216090 800 6 la_data_in[106]
port 125 nsew signal input
rlabel metal2 s 217506 0 217562 800 6 la_data_in[107]
port 126 nsew signal input
rlabel metal2 s 219070 0 219126 800 6 la_data_in[108]
port 127 nsew signal input
rlabel metal2 s 220634 0 220690 800 6 la_data_in[109]
port 128 nsew signal input
rlabel metal2 s 69386 0 69442 800 6 la_data_in[10]
port 129 nsew signal input
rlabel metal2 s 222106 0 222162 800 6 la_data_in[110]
port 130 nsew signal input
rlabel metal2 s 223670 0 223726 800 6 la_data_in[111]
port 131 nsew signal input
rlabel metal2 s 225142 0 225198 800 6 la_data_in[112]
port 132 nsew signal input
rlabel metal2 s 226706 0 226762 800 6 la_data_in[113]
port 133 nsew signal input
rlabel metal2 s 228270 0 228326 800 6 la_data_in[114]
port 134 nsew signal input
rlabel metal2 s 229742 0 229798 800 6 la_data_in[115]
port 135 nsew signal input
rlabel metal2 s 231306 0 231362 800 6 la_data_in[116]
port 136 nsew signal input
rlabel metal2 s 232778 0 232834 800 6 la_data_in[117]
port 137 nsew signal input
rlabel metal2 s 234342 0 234398 800 6 la_data_in[118]
port 138 nsew signal input
rlabel metal2 s 235906 0 235962 800 6 la_data_in[119]
port 139 nsew signal input
rlabel metal2 s 70950 0 71006 800 6 la_data_in[11]
port 140 nsew signal input
rlabel metal2 s 237378 0 237434 800 6 la_data_in[120]
port 141 nsew signal input
rlabel metal2 s 238942 0 238998 800 6 la_data_in[121]
port 142 nsew signal input
rlabel metal2 s 240414 0 240470 800 6 la_data_in[122]
port 143 nsew signal input
rlabel metal2 s 241978 0 242034 800 6 la_data_in[123]
port 144 nsew signal input
rlabel metal2 s 243542 0 243598 800 6 la_data_in[124]
port 145 nsew signal input
rlabel metal2 s 245014 0 245070 800 6 la_data_in[125]
port 146 nsew signal input
rlabel metal2 s 246578 0 246634 800 6 la_data_in[126]
port 147 nsew signal input
rlabel metal2 s 248050 0 248106 800 6 la_data_in[127]
port 148 nsew signal input
rlabel metal2 s 72422 0 72478 800 6 la_data_in[12]
port 149 nsew signal input
rlabel metal2 s 73986 0 74042 800 6 la_data_in[13]
port 150 nsew signal input
rlabel metal2 s 75458 0 75514 800 6 la_data_in[14]
port 151 nsew signal input
rlabel metal2 s 77022 0 77078 800 6 la_data_in[15]
port 152 nsew signal input
rlabel metal2 s 78586 0 78642 800 6 la_data_in[16]
port 153 nsew signal input
rlabel metal2 s 80058 0 80114 800 6 la_data_in[17]
port 154 nsew signal input
rlabel metal2 s 81622 0 81678 800 6 la_data_in[18]
port 155 nsew signal input
rlabel metal2 s 83094 0 83150 800 6 la_data_in[19]
port 156 nsew signal input
rlabel metal2 s 55678 0 55734 800 6 la_data_in[1]
port 157 nsew signal input
rlabel metal2 s 84658 0 84714 800 6 la_data_in[20]
port 158 nsew signal input
rlabel metal2 s 86222 0 86278 800 6 la_data_in[21]
port 159 nsew signal input
rlabel metal2 s 87694 0 87750 800 6 la_data_in[22]
port 160 nsew signal input
rlabel metal2 s 89258 0 89314 800 6 la_data_in[23]
port 161 nsew signal input
rlabel metal2 s 90730 0 90786 800 6 la_data_in[24]
port 162 nsew signal input
rlabel metal2 s 92294 0 92350 800 6 la_data_in[25]
port 163 nsew signal input
rlabel metal2 s 93858 0 93914 800 6 la_data_in[26]
port 164 nsew signal input
rlabel metal2 s 95330 0 95386 800 6 la_data_in[27]
port 165 nsew signal input
rlabel metal2 s 96894 0 96950 800 6 la_data_in[28]
port 166 nsew signal input
rlabel metal2 s 98366 0 98422 800 6 la_data_in[29]
port 167 nsew signal input
rlabel metal2 s 57150 0 57206 800 6 la_data_in[2]
port 168 nsew signal input
rlabel metal2 s 99930 0 99986 800 6 la_data_in[30]
port 169 nsew signal input
rlabel metal2 s 101494 0 101550 800 6 la_data_in[31]
port 170 nsew signal input
rlabel metal2 s 102966 0 103022 800 6 la_data_in[32]
port 171 nsew signal input
rlabel metal2 s 104530 0 104586 800 6 la_data_in[33]
port 172 nsew signal input
rlabel metal2 s 106002 0 106058 800 6 la_data_in[34]
port 173 nsew signal input
rlabel metal2 s 107566 0 107622 800 6 la_data_in[35]
port 174 nsew signal input
rlabel metal2 s 109130 0 109186 800 6 la_data_in[36]
port 175 nsew signal input
rlabel metal2 s 110602 0 110658 800 6 la_data_in[37]
port 176 nsew signal input
rlabel metal2 s 112166 0 112222 800 6 la_data_in[38]
port 177 nsew signal input
rlabel metal2 s 113638 0 113694 800 6 la_data_in[39]
port 178 nsew signal input
rlabel metal2 s 58714 0 58770 800 6 la_data_in[3]
port 179 nsew signal input
rlabel metal2 s 115202 0 115258 800 6 la_data_in[40]
port 180 nsew signal input
rlabel metal2 s 116766 0 116822 800 6 la_data_in[41]
port 181 nsew signal input
rlabel metal2 s 118238 0 118294 800 6 la_data_in[42]
port 182 nsew signal input
rlabel metal2 s 119802 0 119858 800 6 la_data_in[43]
port 183 nsew signal input
rlabel metal2 s 121274 0 121330 800 6 la_data_in[44]
port 184 nsew signal input
rlabel metal2 s 122838 0 122894 800 6 la_data_in[45]
port 185 nsew signal input
rlabel metal2 s 124402 0 124458 800 6 la_data_in[46]
port 186 nsew signal input
rlabel metal2 s 125874 0 125930 800 6 la_data_in[47]
port 187 nsew signal input
rlabel metal2 s 127438 0 127494 800 6 la_data_in[48]
port 188 nsew signal input
rlabel metal2 s 129002 0 129058 800 6 la_data_in[49]
port 189 nsew signal input
rlabel metal2 s 60186 0 60242 800 6 la_data_in[4]
port 190 nsew signal input
rlabel metal2 s 130474 0 130530 800 6 la_data_in[50]
port 191 nsew signal input
rlabel metal2 s 132038 0 132094 800 6 la_data_in[51]
port 192 nsew signal input
rlabel metal2 s 133510 0 133566 800 6 la_data_in[52]
port 193 nsew signal input
rlabel metal2 s 135074 0 135130 800 6 la_data_in[53]
port 194 nsew signal input
rlabel metal2 s 136638 0 136694 800 6 la_data_in[54]
port 195 nsew signal input
rlabel metal2 s 138110 0 138166 800 6 la_data_in[55]
port 196 nsew signal input
rlabel metal2 s 139674 0 139730 800 6 la_data_in[56]
port 197 nsew signal input
rlabel metal2 s 141146 0 141202 800 6 la_data_in[57]
port 198 nsew signal input
rlabel metal2 s 142710 0 142766 800 6 la_data_in[58]
port 199 nsew signal input
rlabel metal2 s 144274 0 144330 800 6 la_data_in[59]
port 200 nsew signal input
rlabel metal2 s 61750 0 61806 800 6 la_data_in[5]
port 201 nsew signal input
rlabel metal2 s 145746 0 145802 800 6 la_data_in[60]
port 202 nsew signal input
rlabel metal2 s 147310 0 147366 800 6 la_data_in[61]
port 203 nsew signal input
rlabel metal2 s 148782 0 148838 800 6 la_data_in[62]
port 204 nsew signal input
rlabel metal2 s 150346 0 150402 800 6 la_data_in[63]
port 205 nsew signal input
rlabel metal2 s 151910 0 151966 800 6 la_data_in[64]
port 206 nsew signal input
rlabel metal2 s 153382 0 153438 800 6 la_data_in[65]
port 207 nsew signal input
rlabel metal2 s 154946 0 155002 800 6 la_data_in[66]
port 208 nsew signal input
rlabel metal2 s 156418 0 156474 800 6 la_data_in[67]
port 209 nsew signal input
rlabel metal2 s 157982 0 158038 800 6 la_data_in[68]
port 210 nsew signal input
rlabel metal2 s 159546 0 159602 800 6 la_data_in[69]
port 211 nsew signal input
rlabel metal2 s 63314 0 63370 800 6 la_data_in[6]
port 212 nsew signal input
rlabel metal2 s 161018 0 161074 800 6 la_data_in[70]
port 213 nsew signal input
rlabel metal2 s 162582 0 162638 800 6 la_data_in[71]
port 214 nsew signal input
rlabel metal2 s 164054 0 164110 800 6 la_data_in[72]
port 215 nsew signal input
rlabel metal2 s 165618 0 165674 800 6 la_data_in[73]
port 216 nsew signal input
rlabel metal2 s 167182 0 167238 800 6 la_data_in[74]
port 217 nsew signal input
rlabel metal2 s 168654 0 168710 800 6 la_data_in[75]
port 218 nsew signal input
rlabel metal2 s 170218 0 170274 800 6 la_data_in[76]
port 219 nsew signal input
rlabel metal2 s 171690 0 171746 800 6 la_data_in[77]
port 220 nsew signal input
rlabel metal2 s 173254 0 173310 800 6 la_data_in[78]
port 221 nsew signal input
rlabel metal2 s 174818 0 174874 800 6 la_data_in[79]
port 222 nsew signal input
rlabel metal2 s 64786 0 64842 800 6 la_data_in[7]
port 223 nsew signal input
rlabel metal2 s 176290 0 176346 800 6 la_data_in[80]
port 224 nsew signal input
rlabel metal2 s 177854 0 177910 800 6 la_data_in[81]
port 225 nsew signal input
rlabel metal2 s 179326 0 179382 800 6 la_data_in[82]
port 226 nsew signal input
rlabel metal2 s 180890 0 180946 800 6 la_data_in[83]
port 227 nsew signal input
rlabel metal2 s 182454 0 182510 800 6 la_data_in[84]
port 228 nsew signal input
rlabel metal2 s 183926 0 183982 800 6 la_data_in[85]
port 229 nsew signal input
rlabel metal2 s 185490 0 185546 800 6 la_data_in[86]
port 230 nsew signal input
rlabel metal2 s 186962 0 187018 800 6 la_data_in[87]
port 231 nsew signal input
rlabel metal2 s 188526 0 188582 800 6 la_data_in[88]
port 232 nsew signal input
rlabel metal2 s 190090 0 190146 800 6 la_data_in[89]
port 233 nsew signal input
rlabel metal2 s 66350 0 66406 800 6 la_data_in[8]
port 234 nsew signal input
rlabel metal2 s 191562 0 191618 800 6 la_data_in[90]
port 235 nsew signal input
rlabel metal2 s 193126 0 193182 800 6 la_data_in[91]
port 236 nsew signal input
rlabel metal2 s 194598 0 194654 800 6 la_data_in[92]
port 237 nsew signal input
rlabel metal2 s 196162 0 196218 800 6 la_data_in[93]
port 238 nsew signal input
rlabel metal2 s 197726 0 197782 800 6 la_data_in[94]
port 239 nsew signal input
rlabel metal2 s 199198 0 199254 800 6 la_data_in[95]
port 240 nsew signal input
rlabel metal2 s 200762 0 200818 800 6 la_data_in[96]
port 241 nsew signal input
rlabel metal2 s 202234 0 202290 800 6 la_data_in[97]
port 242 nsew signal input
rlabel metal2 s 203798 0 203854 800 6 la_data_in[98]
port 243 nsew signal input
rlabel metal2 s 205362 0 205418 800 6 la_data_in[99]
port 244 nsew signal input
rlabel metal2 s 67822 0 67878 800 6 la_data_in[9]
port 245 nsew signal input
rlabel metal2 s 54666 0 54722 800 6 la_data_out[0]
port 246 nsew signal output
rlabel metal2 s 207386 0 207442 800 6 la_data_out[100]
port 247 nsew signal output
rlabel metal2 s 208858 0 208914 800 6 la_data_out[101]
port 248 nsew signal output
rlabel metal2 s 210422 0 210478 800 6 la_data_out[102]
port 249 nsew signal output
rlabel metal2 s 211894 0 211950 800 6 la_data_out[103]
port 250 nsew signal output
rlabel metal2 s 213458 0 213514 800 6 la_data_out[104]
port 251 nsew signal output
rlabel metal2 s 215022 0 215078 800 6 la_data_out[105]
port 252 nsew signal output
rlabel metal2 s 216494 0 216550 800 6 la_data_out[106]
port 253 nsew signal output
rlabel metal2 s 218058 0 218114 800 6 la_data_out[107]
port 254 nsew signal output
rlabel metal2 s 219530 0 219586 800 6 la_data_out[108]
port 255 nsew signal output
rlabel metal2 s 221094 0 221150 800 6 la_data_out[109]
port 256 nsew signal output
rlabel metal2 s 69938 0 69994 800 6 la_data_out[10]
port 257 nsew signal output
rlabel metal2 s 222658 0 222714 800 6 la_data_out[110]
port 258 nsew signal output
rlabel metal2 s 224130 0 224186 800 6 la_data_out[111]
port 259 nsew signal output
rlabel metal2 s 225694 0 225750 800 6 la_data_out[112]
port 260 nsew signal output
rlabel metal2 s 227166 0 227222 800 6 la_data_out[113]
port 261 nsew signal output
rlabel metal2 s 228730 0 228786 800 6 la_data_out[114]
port 262 nsew signal output
rlabel metal2 s 230294 0 230350 800 6 la_data_out[115]
port 263 nsew signal output
rlabel metal2 s 231766 0 231822 800 6 la_data_out[116]
port 264 nsew signal output
rlabel metal2 s 233330 0 233386 800 6 la_data_out[117]
port 265 nsew signal output
rlabel metal2 s 234802 0 234858 800 6 la_data_out[118]
port 266 nsew signal output
rlabel metal2 s 236366 0 236422 800 6 la_data_out[119]
port 267 nsew signal output
rlabel metal2 s 71410 0 71466 800 6 la_data_out[11]
port 268 nsew signal output
rlabel metal2 s 237930 0 237986 800 6 la_data_out[120]
port 269 nsew signal output
rlabel metal2 s 239402 0 239458 800 6 la_data_out[121]
port 270 nsew signal output
rlabel metal2 s 240966 0 241022 800 6 la_data_out[122]
port 271 nsew signal output
rlabel metal2 s 242438 0 242494 800 6 la_data_out[123]
port 272 nsew signal output
rlabel metal2 s 244002 0 244058 800 6 la_data_out[124]
port 273 nsew signal output
rlabel metal2 s 245566 0 245622 800 6 la_data_out[125]
port 274 nsew signal output
rlabel metal2 s 247038 0 247094 800 6 la_data_out[126]
port 275 nsew signal output
rlabel metal2 s 248602 0 248658 800 6 la_data_out[127]
port 276 nsew signal output
rlabel metal2 s 72974 0 73030 800 6 la_data_out[12]
port 277 nsew signal output
rlabel metal2 s 74446 0 74502 800 6 la_data_out[13]
port 278 nsew signal output
rlabel metal2 s 76010 0 76066 800 6 la_data_out[14]
port 279 nsew signal output
rlabel metal2 s 77574 0 77630 800 6 la_data_out[15]
port 280 nsew signal output
rlabel metal2 s 79046 0 79102 800 6 la_data_out[16]
port 281 nsew signal output
rlabel metal2 s 80610 0 80666 800 6 la_data_out[17]
port 282 nsew signal output
rlabel metal2 s 82082 0 82138 800 6 la_data_out[18]
port 283 nsew signal output
rlabel metal2 s 83646 0 83702 800 6 la_data_out[19]
port 284 nsew signal output
rlabel metal2 s 56138 0 56194 800 6 la_data_out[1]
port 285 nsew signal output
rlabel metal2 s 85210 0 85266 800 6 la_data_out[20]
port 286 nsew signal output
rlabel metal2 s 86682 0 86738 800 6 la_data_out[21]
port 287 nsew signal output
rlabel metal2 s 88246 0 88302 800 6 la_data_out[22]
port 288 nsew signal output
rlabel metal2 s 89718 0 89774 800 6 la_data_out[23]
port 289 nsew signal output
rlabel metal2 s 91282 0 91338 800 6 la_data_out[24]
port 290 nsew signal output
rlabel metal2 s 92846 0 92902 800 6 la_data_out[25]
port 291 nsew signal output
rlabel metal2 s 94318 0 94374 800 6 la_data_out[26]
port 292 nsew signal output
rlabel metal2 s 95882 0 95938 800 6 la_data_out[27]
port 293 nsew signal output
rlabel metal2 s 97354 0 97410 800 6 la_data_out[28]
port 294 nsew signal output
rlabel metal2 s 98918 0 98974 800 6 la_data_out[29]
port 295 nsew signal output
rlabel metal2 s 57702 0 57758 800 6 la_data_out[2]
port 296 nsew signal output
rlabel metal2 s 100482 0 100538 800 6 la_data_out[30]
port 297 nsew signal output
rlabel metal2 s 101954 0 102010 800 6 la_data_out[31]
port 298 nsew signal output
rlabel metal2 s 103518 0 103574 800 6 la_data_out[32]
port 299 nsew signal output
rlabel metal2 s 104990 0 105046 800 6 la_data_out[33]
port 300 nsew signal output
rlabel metal2 s 106554 0 106610 800 6 la_data_out[34]
port 301 nsew signal output
rlabel metal2 s 108118 0 108174 800 6 la_data_out[35]
port 302 nsew signal output
rlabel metal2 s 109590 0 109646 800 6 la_data_out[36]
port 303 nsew signal output
rlabel metal2 s 111154 0 111210 800 6 la_data_out[37]
port 304 nsew signal output
rlabel metal2 s 112626 0 112682 800 6 la_data_out[38]
port 305 nsew signal output
rlabel metal2 s 114190 0 114246 800 6 la_data_out[39]
port 306 nsew signal output
rlabel metal2 s 59174 0 59230 800 6 la_data_out[3]
port 307 nsew signal output
rlabel metal2 s 115754 0 115810 800 6 la_data_out[40]
port 308 nsew signal output
rlabel metal2 s 117226 0 117282 800 6 la_data_out[41]
port 309 nsew signal output
rlabel metal2 s 118790 0 118846 800 6 la_data_out[42]
port 310 nsew signal output
rlabel metal2 s 120262 0 120318 800 6 la_data_out[43]
port 311 nsew signal output
rlabel metal2 s 121826 0 121882 800 6 la_data_out[44]
port 312 nsew signal output
rlabel metal2 s 123390 0 123446 800 6 la_data_out[45]
port 313 nsew signal output
rlabel metal2 s 124862 0 124918 800 6 la_data_out[46]
port 314 nsew signal output
rlabel metal2 s 126426 0 126482 800 6 la_data_out[47]
port 315 nsew signal output
rlabel metal2 s 127898 0 127954 800 6 la_data_out[48]
port 316 nsew signal output
rlabel metal2 s 129462 0 129518 800 6 la_data_out[49]
port 317 nsew signal output
rlabel metal2 s 60738 0 60794 800 6 la_data_out[4]
port 318 nsew signal output
rlabel metal2 s 131026 0 131082 800 6 la_data_out[50]
port 319 nsew signal output
rlabel metal2 s 132498 0 132554 800 6 la_data_out[51]
port 320 nsew signal output
rlabel metal2 s 134062 0 134118 800 6 la_data_out[52]
port 321 nsew signal output
rlabel metal2 s 135534 0 135590 800 6 la_data_out[53]
port 322 nsew signal output
rlabel metal2 s 137098 0 137154 800 6 la_data_out[54]
port 323 nsew signal output
rlabel metal2 s 138662 0 138718 800 6 la_data_out[55]
port 324 nsew signal output
rlabel metal2 s 140134 0 140190 800 6 la_data_out[56]
port 325 nsew signal output
rlabel metal2 s 141698 0 141754 800 6 la_data_out[57]
port 326 nsew signal output
rlabel metal2 s 143170 0 143226 800 6 la_data_out[58]
port 327 nsew signal output
rlabel metal2 s 144734 0 144790 800 6 la_data_out[59]
port 328 nsew signal output
rlabel metal2 s 62302 0 62358 800 6 la_data_out[5]
port 329 nsew signal output
rlabel metal2 s 146298 0 146354 800 6 la_data_out[60]
port 330 nsew signal output
rlabel metal2 s 147770 0 147826 800 6 la_data_out[61]
port 331 nsew signal output
rlabel metal2 s 149334 0 149390 800 6 la_data_out[62]
port 332 nsew signal output
rlabel metal2 s 150806 0 150862 800 6 la_data_out[63]
port 333 nsew signal output
rlabel metal2 s 152370 0 152426 800 6 la_data_out[64]
port 334 nsew signal output
rlabel metal2 s 153934 0 153990 800 6 la_data_out[65]
port 335 nsew signal output
rlabel metal2 s 155406 0 155462 800 6 la_data_out[66]
port 336 nsew signal output
rlabel metal2 s 156970 0 157026 800 6 la_data_out[67]
port 337 nsew signal output
rlabel metal2 s 158442 0 158498 800 6 la_data_out[68]
port 338 nsew signal output
rlabel metal2 s 160006 0 160062 800 6 la_data_out[69]
port 339 nsew signal output
rlabel metal2 s 63774 0 63830 800 6 la_data_out[6]
port 340 nsew signal output
rlabel metal2 s 161570 0 161626 800 6 la_data_out[70]
port 341 nsew signal output
rlabel metal2 s 163042 0 163098 800 6 la_data_out[71]
port 342 nsew signal output
rlabel metal2 s 164606 0 164662 800 6 la_data_out[72]
port 343 nsew signal output
rlabel metal2 s 166078 0 166134 800 6 la_data_out[73]
port 344 nsew signal output
rlabel metal2 s 167642 0 167698 800 6 la_data_out[74]
port 345 nsew signal output
rlabel metal2 s 169206 0 169262 800 6 la_data_out[75]
port 346 nsew signal output
rlabel metal2 s 170678 0 170734 800 6 la_data_out[76]
port 347 nsew signal output
rlabel metal2 s 172242 0 172298 800 6 la_data_out[77]
port 348 nsew signal output
rlabel metal2 s 173714 0 173770 800 6 la_data_out[78]
port 349 nsew signal output
rlabel metal2 s 175278 0 175334 800 6 la_data_out[79]
port 350 nsew signal output
rlabel metal2 s 65338 0 65394 800 6 la_data_out[7]
port 351 nsew signal output
rlabel metal2 s 176842 0 176898 800 6 la_data_out[80]
port 352 nsew signal output
rlabel metal2 s 178314 0 178370 800 6 la_data_out[81]
port 353 nsew signal output
rlabel metal2 s 179878 0 179934 800 6 la_data_out[82]
port 354 nsew signal output
rlabel metal2 s 181350 0 181406 800 6 la_data_out[83]
port 355 nsew signal output
rlabel metal2 s 182914 0 182970 800 6 la_data_out[84]
port 356 nsew signal output
rlabel metal2 s 184478 0 184534 800 6 la_data_out[85]
port 357 nsew signal output
rlabel metal2 s 185950 0 186006 800 6 la_data_out[86]
port 358 nsew signal output
rlabel metal2 s 187514 0 187570 800 6 la_data_out[87]
port 359 nsew signal output
rlabel metal2 s 188986 0 189042 800 6 la_data_out[88]
port 360 nsew signal output
rlabel metal2 s 190550 0 190606 800 6 la_data_out[89]
port 361 nsew signal output
rlabel metal2 s 66810 0 66866 800 6 la_data_out[8]
port 362 nsew signal output
rlabel metal2 s 192114 0 192170 800 6 la_data_out[90]
port 363 nsew signal output
rlabel metal2 s 193586 0 193642 800 6 la_data_out[91]
port 364 nsew signal output
rlabel metal2 s 195150 0 195206 800 6 la_data_out[92]
port 365 nsew signal output
rlabel metal2 s 196622 0 196678 800 6 la_data_out[93]
port 366 nsew signal output
rlabel metal2 s 198186 0 198242 800 6 la_data_out[94]
port 367 nsew signal output
rlabel metal2 s 199750 0 199806 800 6 la_data_out[95]
port 368 nsew signal output
rlabel metal2 s 201222 0 201278 800 6 la_data_out[96]
port 369 nsew signal output
rlabel metal2 s 202786 0 202842 800 6 la_data_out[97]
port 370 nsew signal output
rlabel metal2 s 204258 0 204314 800 6 la_data_out[98]
port 371 nsew signal output
rlabel metal2 s 205822 0 205878 800 6 la_data_out[99]
port 372 nsew signal output
rlabel metal2 s 68374 0 68430 800 6 la_data_out[9]
port 373 nsew signal output
rlabel metal2 s 55126 0 55182 800 6 la_oenb[0]
port 374 nsew signal input
rlabel metal2 s 207846 0 207902 800 6 la_oenb[100]
port 375 nsew signal input
rlabel metal2 s 209410 0 209466 800 6 la_oenb[101]
port 376 nsew signal input
rlabel metal2 s 210882 0 210938 800 6 la_oenb[102]
port 377 nsew signal input
rlabel metal2 s 212446 0 212502 800 6 la_oenb[103]
port 378 nsew signal input
rlabel metal2 s 214010 0 214066 800 6 la_oenb[104]
port 379 nsew signal input
rlabel metal2 s 215482 0 215538 800 6 la_oenb[105]
port 380 nsew signal input
rlabel metal2 s 217046 0 217102 800 6 la_oenb[106]
port 381 nsew signal input
rlabel metal2 s 218518 0 218574 800 6 la_oenb[107]
port 382 nsew signal input
rlabel metal2 s 220082 0 220138 800 6 la_oenb[108]
port 383 nsew signal input
rlabel metal2 s 221646 0 221702 800 6 la_oenb[109]
port 384 nsew signal input
rlabel metal2 s 70398 0 70454 800 6 la_oenb[10]
port 385 nsew signal input
rlabel metal2 s 223118 0 223174 800 6 la_oenb[110]
port 386 nsew signal input
rlabel metal2 s 224682 0 224738 800 6 la_oenb[111]
port 387 nsew signal input
rlabel metal2 s 226154 0 226210 800 6 la_oenb[112]
port 388 nsew signal input
rlabel metal2 s 227718 0 227774 800 6 la_oenb[113]
port 389 nsew signal input
rlabel metal2 s 229282 0 229338 800 6 la_oenb[114]
port 390 nsew signal input
rlabel metal2 s 230754 0 230810 800 6 la_oenb[115]
port 391 nsew signal input
rlabel metal2 s 232318 0 232374 800 6 la_oenb[116]
port 392 nsew signal input
rlabel metal2 s 233790 0 233846 800 6 la_oenb[117]
port 393 nsew signal input
rlabel metal2 s 235354 0 235410 800 6 la_oenb[118]
port 394 nsew signal input
rlabel metal2 s 236918 0 236974 800 6 la_oenb[119]
port 395 nsew signal input
rlabel metal2 s 71962 0 72018 800 6 la_oenb[11]
port 396 nsew signal input
rlabel metal2 s 238390 0 238446 800 6 la_oenb[120]
port 397 nsew signal input
rlabel metal2 s 239954 0 240010 800 6 la_oenb[121]
port 398 nsew signal input
rlabel metal2 s 241426 0 241482 800 6 la_oenb[122]
port 399 nsew signal input
rlabel metal2 s 242990 0 243046 800 6 la_oenb[123]
port 400 nsew signal input
rlabel metal2 s 244554 0 244610 800 6 la_oenb[124]
port 401 nsew signal input
rlabel metal2 s 246026 0 246082 800 6 la_oenb[125]
port 402 nsew signal input
rlabel metal2 s 247590 0 247646 800 6 la_oenb[126]
port 403 nsew signal input
rlabel metal2 s 249062 0 249118 800 6 la_oenb[127]
port 404 nsew signal input
rlabel metal2 s 73434 0 73490 800 6 la_oenb[12]
port 405 nsew signal input
rlabel metal2 s 74998 0 75054 800 6 la_oenb[13]
port 406 nsew signal input
rlabel metal2 s 76562 0 76618 800 6 la_oenb[14]
port 407 nsew signal input
rlabel metal2 s 78034 0 78090 800 6 la_oenb[15]
port 408 nsew signal input
rlabel metal2 s 79598 0 79654 800 6 la_oenb[16]
port 409 nsew signal input
rlabel metal2 s 81070 0 81126 800 6 la_oenb[17]
port 410 nsew signal input
rlabel metal2 s 82634 0 82690 800 6 la_oenb[18]
port 411 nsew signal input
rlabel metal2 s 84198 0 84254 800 6 la_oenb[19]
port 412 nsew signal input
rlabel metal2 s 56690 0 56746 800 6 la_oenb[1]
port 413 nsew signal input
rlabel metal2 s 85670 0 85726 800 6 la_oenb[20]
port 414 nsew signal input
rlabel metal2 s 87234 0 87290 800 6 la_oenb[21]
port 415 nsew signal input
rlabel metal2 s 88706 0 88762 800 6 la_oenb[22]
port 416 nsew signal input
rlabel metal2 s 90270 0 90326 800 6 la_oenb[23]
port 417 nsew signal input
rlabel metal2 s 91834 0 91890 800 6 la_oenb[24]
port 418 nsew signal input
rlabel metal2 s 93306 0 93362 800 6 la_oenb[25]
port 419 nsew signal input
rlabel metal2 s 94870 0 94926 800 6 la_oenb[26]
port 420 nsew signal input
rlabel metal2 s 96342 0 96398 800 6 la_oenb[27]
port 421 nsew signal input
rlabel metal2 s 97906 0 97962 800 6 la_oenb[28]
port 422 nsew signal input
rlabel metal2 s 99470 0 99526 800 6 la_oenb[29]
port 423 nsew signal input
rlabel metal2 s 58162 0 58218 800 6 la_oenb[2]
port 424 nsew signal input
rlabel metal2 s 100942 0 100998 800 6 la_oenb[30]
port 425 nsew signal input
rlabel metal2 s 102506 0 102562 800 6 la_oenb[31]
port 426 nsew signal input
rlabel metal2 s 103978 0 104034 800 6 la_oenb[32]
port 427 nsew signal input
rlabel metal2 s 105542 0 105598 800 6 la_oenb[33]
port 428 nsew signal input
rlabel metal2 s 107106 0 107162 800 6 la_oenb[34]
port 429 nsew signal input
rlabel metal2 s 108578 0 108634 800 6 la_oenb[35]
port 430 nsew signal input
rlabel metal2 s 110142 0 110198 800 6 la_oenb[36]
port 431 nsew signal input
rlabel metal2 s 111614 0 111670 800 6 la_oenb[37]
port 432 nsew signal input
rlabel metal2 s 113178 0 113234 800 6 la_oenb[38]
port 433 nsew signal input
rlabel metal2 s 114742 0 114798 800 6 la_oenb[39]
port 434 nsew signal input
rlabel metal2 s 59726 0 59782 800 6 la_oenb[3]
port 435 nsew signal input
rlabel metal2 s 116214 0 116270 800 6 la_oenb[40]
port 436 nsew signal input
rlabel metal2 s 117778 0 117834 800 6 la_oenb[41]
port 437 nsew signal input
rlabel metal2 s 119250 0 119306 800 6 la_oenb[42]
port 438 nsew signal input
rlabel metal2 s 120814 0 120870 800 6 la_oenb[43]
port 439 nsew signal input
rlabel metal2 s 122378 0 122434 800 6 la_oenb[44]
port 440 nsew signal input
rlabel metal2 s 123850 0 123906 800 6 la_oenb[45]
port 441 nsew signal input
rlabel metal2 s 125414 0 125470 800 6 la_oenb[46]
port 442 nsew signal input
rlabel metal2 s 126886 0 126942 800 6 la_oenb[47]
port 443 nsew signal input
rlabel metal2 s 128450 0 128506 800 6 la_oenb[48]
port 444 nsew signal input
rlabel metal2 s 130014 0 130070 800 6 la_oenb[49]
port 445 nsew signal input
rlabel metal2 s 61290 0 61346 800 6 la_oenb[4]
port 446 nsew signal input
rlabel metal2 s 131486 0 131542 800 6 la_oenb[50]
port 447 nsew signal input
rlabel metal2 s 133050 0 133106 800 6 la_oenb[51]
port 448 nsew signal input
rlabel metal2 s 134522 0 134578 800 6 la_oenb[52]
port 449 nsew signal input
rlabel metal2 s 136086 0 136142 800 6 la_oenb[53]
port 450 nsew signal input
rlabel metal2 s 137650 0 137706 800 6 la_oenb[54]
port 451 nsew signal input
rlabel metal2 s 139122 0 139178 800 6 la_oenb[55]
port 452 nsew signal input
rlabel metal2 s 140686 0 140742 800 6 la_oenb[56]
port 453 nsew signal input
rlabel metal2 s 142158 0 142214 800 6 la_oenb[57]
port 454 nsew signal input
rlabel metal2 s 143722 0 143778 800 6 la_oenb[58]
port 455 nsew signal input
rlabel metal2 s 145286 0 145342 800 6 la_oenb[59]
port 456 nsew signal input
rlabel metal2 s 62762 0 62818 800 6 la_oenb[5]
port 457 nsew signal input
rlabel metal2 s 146758 0 146814 800 6 la_oenb[60]
port 458 nsew signal input
rlabel metal2 s 148322 0 148378 800 6 la_oenb[61]
port 459 nsew signal input
rlabel metal2 s 149794 0 149850 800 6 la_oenb[62]
port 460 nsew signal input
rlabel metal2 s 151358 0 151414 800 6 la_oenb[63]
port 461 nsew signal input
rlabel metal2 s 152922 0 152978 800 6 la_oenb[64]
port 462 nsew signal input
rlabel metal2 s 154394 0 154450 800 6 la_oenb[65]
port 463 nsew signal input
rlabel metal2 s 155958 0 156014 800 6 la_oenb[66]
port 464 nsew signal input
rlabel metal2 s 157430 0 157486 800 6 la_oenb[67]
port 465 nsew signal input
rlabel metal2 s 158994 0 159050 800 6 la_oenb[68]
port 466 nsew signal input
rlabel metal2 s 160558 0 160614 800 6 la_oenb[69]
port 467 nsew signal input
rlabel metal2 s 64326 0 64382 800 6 la_oenb[6]
port 468 nsew signal input
rlabel metal2 s 162030 0 162086 800 6 la_oenb[70]
port 469 nsew signal input
rlabel metal2 s 163594 0 163650 800 6 la_oenb[71]
port 470 nsew signal input
rlabel metal2 s 165066 0 165122 800 6 la_oenb[72]
port 471 nsew signal input
rlabel metal2 s 166630 0 166686 800 6 la_oenb[73]
port 472 nsew signal input
rlabel metal2 s 168194 0 168250 800 6 la_oenb[74]
port 473 nsew signal input
rlabel metal2 s 169666 0 169722 800 6 la_oenb[75]
port 474 nsew signal input
rlabel metal2 s 171230 0 171286 800 6 la_oenb[76]
port 475 nsew signal input
rlabel metal2 s 172702 0 172758 800 6 la_oenb[77]
port 476 nsew signal input
rlabel metal2 s 174266 0 174322 800 6 la_oenb[78]
port 477 nsew signal input
rlabel metal2 s 175830 0 175886 800 6 la_oenb[79]
port 478 nsew signal input
rlabel metal2 s 65798 0 65854 800 6 la_oenb[7]
port 479 nsew signal input
rlabel metal2 s 177302 0 177358 800 6 la_oenb[80]
port 480 nsew signal input
rlabel metal2 s 178866 0 178922 800 6 la_oenb[81]
port 481 nsew signal input
rlabel metal2 s 180338 0 180394 800 6 la_oenb[82]
port 482 nsew signal input
rlabel metal2 s 181902 0 181958 800 6 la_oenb[83]
port 483 nsew signal input
rlabel metal2 s 183466 0 183522 800 6 la_oenb[84]
port 484 nsew signal input
rlabel metal2 s 184938 0 184994 800 6 la_oenb[85]
port 485 nsew signal input
rlabel metal2 s 186502 0 186558 800 6 la_oenb[86]
port 486 nsew signal input
rlabel metal2 s 187974 0 188030 800 6 la_oenb[87]
port 487 nsew signal input
rlabel metal2 s 189538 0 189594 800 6 la_oenb[88]
port 488 nsew signal input
rlabel metal2 s 191102 0 191158 800 6 la_oenb[89]
port 489 nsew signal input
rlabel metal2 s 67362 0 67418 800 6 la_oenb[8]
port 490 nsew signal input
rlabel metal2 s 192574 0 192630 800 6 la_oenb[90]
port 491 nsew signal input
rlabel metal2 s 194138 0 194194 800 6 la_oenb[91]
port 492 nsew signal input
rlabel metal2 s 195610 0 195666 800 6 la_oenb[92]
port 493 nsew signal input
rlabel metal2 s 197174 0 197230 800 6 la_oenb[93]
port 494 nsew signal input
rlabel metal2 s 198738 0 198794 800 6 la_oenb[94]
port 495 nsew signal input
rlabel metal2 s 200210 0 200266 800 6 la_oenb[95]
port 496 nsew signal input
rlabel metal2 s 201774 0 201830 800 6 la_oenb[96]
port 497 nsew signal input
rlabel metal2 s 203246 0 203302 800 6 la_oenb[97]
port 498 nsew signal input
rlabel metal2 s 204810 0 204866 800 6 la_oenb[98]
port 499 nsew signal input
rlabel metal2 s 206374 0 206430 800 6 la_oenb[99]
port 500 nsew signal input
rlabel metal2 s 68926 0 68982 800 6 la_oenb[9]
port 501 nsew signal input
rlabel metal4 s 4208 2128 4528 247568 6 vccd1
port 502 nsew power input
rlabel metal4 s 34928 2128 35248 247568 6 vccd1
port 502 nsew power input
rlabel metal4 s 65648 2128 65968 247568 6 vccd1
port 502 nsew power input
rlabel metal4 s 96368 2128 96688 247568 6 vccd1
port 502 nsew power input
rlabel metal4 s 127088 2128 127408 247568 6 vccd1
port 502 nsew power input
rlabel metal4 s 157808 2128 158128 247568 6 vccd1
port 502 nsew power input
rlabel metal4 s 188528 2128 188848 247568 6 vccd1
port 502 nsew power input
rlabel metal4 s 219248 2128 219568 247568 6 vccd1
port 502 nsew power input
rlabel metal4 s 19568 2128 19888 247568 6 vssd1
port 503 nsew ground input
rlabel metal4 s 50288 2128 50608 247568 6 vssd1
port 503 nsew ground input
rlabel metal4 s 81008 2128 81328 247568 6 vssd1
port 503 nsew ground input
rlabel metal4 s 111728 2128 112048 247568 6 vssd1
port 503 nsew ground input
rlabel metal4 s 142448 2128 142768 247568 6 vssd1
port 503 nsew ground input
rlabel metal4 s 173168 2128 173488 247568 6 vssd1
port 503 nsew ground input
rlabel metal4 s 203888 2128 204208 247568 6 vssd1
port 503 nsew ground input
rlabel metal4 s 234608 2128 234928 247568 6 vssd1
port 503 nsew ground input
rlabel metal2 s 202 0 258 800 6 wb_clk_i
port 504 nsew signal input
rlabel metal2 s 662 0 718 800 6 wb_rst_i
port 505 nsew signal input
rlabel metal2 s 1214 0 1270 800 6 wbs_ack_o
port 506 nsew signal output
rlabel metal2 s 3238 0 3294 800 6 wbs_adr_i[0]
port 507 nsew signal input
rlabel metal2 s 20534 0 20590 800 6 wbs_adr_i[10]
port 508 nsew signal input
rlabel metal2 s 22006 0 22062 800 6 wbs_adr_i[11]
port 509 nsew signal input
rlabel metal2 s 23570 0 23626 800 6 wbs_adr_i[12]
port 510 nsew signal input
rlabel metal2 s 25134 0 25190 800 6 wbs_adr_i[13]
port 511 nsew signal input
rlabel metal2 s 26606 0 26662 800 6 wbs_adr_i[14]
port 512 nsew signal input
rlabel metal2 s 28170 0 28226 800 6 wbs_adr_i[15]
port 513 nsew signal input
rlabel metal2 s 29642 0 29698 800 6 wbs_adr_i[16]
port 514 nsew signal input
rlabel metal2 s 31206 0 31262 800 6 wbs_adr_i[17]
port 515 nsew signal input
rlabel metal2 s 32770 0 32826 800 6 wbs_adr_i[18]
port 516 nsew signal input
rlabel metal2 s 34242 0 34298 800 6 wbs_adr_i[19]
port 517 nsew signal input
rlabel metal2 s 5262 0 5318 800 6 wbs_adr_i[1]
port 518 nsew signal input
rlabel metal2 s 35806 0 35862 800 6 wbs_adr_i[20]
port 519 nsew signal input
rlabel metal2 s 37278 0 37334 800 6 wbs_adr_i[21]
port 520 nsew signal input
rlabel metal2 s 38842 0 38898 800 6 wbs_adr_i[22]
port 521 nsew signal input
rlabel metal2 s 40406 0 40462 800 6 wbs_adr_i[23]
port 522 nsew signal input
rlabel metal2 s 41878 0 41934 800 6 wbs_adr_i[24]
port 523 nsew signal input
rlabel metal2 s 43442 0 43498 800 6 wbs_adr_i[25]
port 524 nsew signal input
rlabel metal2 s 44914 0 44970 800 6 wbs_adr_i[26]
port 525 nsew signal input
rlabel metal2 s 46478 0 46534 800 6 wbs_adr_i[27]
port 526 nsew signal input
rlabel metal2 s 48042 0 48098 800 6 wbs_adr_i[28]
port 527 nsew signal input
rlabel metal2 s 49514 0 49570 800 6 wbs_adr_i[29]
port 528 nsew signal input
rlabel metal2 s 7286 0 7342 800 6 wbs_adr_i[2]
port 529 nsew signal input
rlabel metal2 s 51078 0 51134 800 6 wbs_adr_i[30]
port 530 nsew signal input
rlabel metal2 s 52550 0 52606 800 6 wbs_adr_i[31]
port 531 nsew signal input
rlabel metal2 s 9310 0 9366 800 6 wbs_adr_i[3]
port 532 nsew signal input
rlabel metal2 s 11334 0 11390 800 6 wbs_adr_i[4]
port 533 nsew signal input
rlabel metal2 s 12898 0 12954 800 6 wbs_adr_i[5]
port 534 nsew signal input
rlabel metal2 s 14370 0 14426 800 6 wbs_adr_i[6]
port 535 nsew signal input
rlabel metal2 s 15934 0 15990 800 6 wbs_adr_i[7]
port 536 nsew signal input
rlabel metal2 s 17498 0 17554 800 6 wbs_adr_i[8]
port 537 nsew signal input
rlabel metal2 s 18970 0 19026 800 6 wbs_adr_i[9]
port 538 nsew signal input
rlabel metal2 s 1674 0 1730 800 6 wbs_cyc_i
port 539 nsew signal input
rlabel metal2 s 3698 0 3754 800 6 wbs_dat_i[0]
port 540 nsew signal input
rlabel metal2 s 20994 0 21050 800 6 wbs_dat_i[10]
port 541 nsew signal input
rlabel metal2 s 22558 0 22614 800 6 wbs_dat_i[11]
port 542 nsew signal input
rlabel metal2 s 24122 0 24178 800 6 wbs_dat_i[12]
port 543 nsew signal input
rlabel metal2 s 25594 0 25650 800 6 wbs_dat_i[13]
port 544 nsew signal input
rlabel metal2 s 27158 0 27214 800 6 wbs_dat_i[14]
port 545 nsew signal input
rlabel metal2 s 28630 0 28686 800 6 wbs_dat_i[15]
port 546 nsew signal input
rlabel metal2 s 30194 0 30250 800 6 wbs_dat_i[16]
port 547 nsew signal input
rlabel metal2 s 31758 0 31814 800 6 wbs_dat_i[17]
port 548 nsew signal input
rlabel metal2 s 33230 0 33286 800 6 wbs_dat_i[18]
port 549 nsew signal input
rlabel metal2 s 34794 0 34850 800 6 wbs_dat_i[19]
port 550 nsew signal input
rlabel metal2 s 5722 0 5778 800 6 wbs_dat_i[1]
port 551 nsew signal input
rlabel metal2 s 36266 0 36322 800 6 wbs_dat_i[20]
port 552 nsew signal input
rlabel metal2 s 37830 0 37886 800 6 wbs_dat_i[21]
port 553 nsew signal input
rlabel metal2 s 39394 0 39450 800 6 wbs_dat_i[22]
port 554 nsew signal input
rlabel metal2 s 40866 0 40922 800 6 wbs_dat_i[23]
port 555 nsew signal input
rlabel metal2 s 42430 0 42486 800 6 wbs_dat_i[24]
port 556 nsew signal input
rlabel metal2 s 43902 0 43958 800 6 wbs_dat_i[25]
port 557 nsew signal input
rlabel metal2 s 45466 0 45522 800 6 wbs_dat_i[26]
port 558 nsew signal input
rlabel metal2 s 47030 0 47086 800 6 wbs_dat_i[27]
port 559 nsew signal input
rlabel metal2 s 48502 0 48558 800 6 wbs_dat_i[28]
port 560 nsew signal input
rlabel metal2 s 50066 0 50122 800 6 wbs_dat_i[29]
port 561 nsew signal input
rlabel metal2 s 7838 0 7894 800 6 wbs_dat_i[2]
port 562 nsew signal input
rlabel metal2 s 51538 0 51594 800 6 wbs_dat_i[30]
port 563 nsew signal input
rlabel metal2 s 53102 0 53158 800 6 wbs_dat_i[31]
port 564 nsew signal input
rlabel metal2 s 9862 0 9918 800 6 wbs_dat_i[3]
port 565 nsew signal input
rlabel metal2 s 11886 0 11942 800 6 wbs_dat_i[4]
port 566 nsew signal input
rlabel metal2 s 13358 0 13414 800 6 wbs_dat_i[5]
port 567 nsew signal input
rlabel metal2 s 14922 0 14978 800 6 wbs_dat_i[6]
port 568 nsew signal input
rlabel metal2 s 16486 0 16542 800 6 wbs_dat_i[7]
port 569 nsew signal input
rlabel metal2 s 17958 0 18014 800 6 wbs_dat_i[8]
port 570 nsew signal input
rlabel metal2 s 19522 0 19578 800 6 wbs_dat_i[9]
port 571 nsew signal input
rlabel metal2 s 4250 0 4306 800 6 wbs_dat_o[0]
port 572 nsew signal output
rlabel metal2 s 21546 0 21602 800 6 wbs_dat_o[10]
port 573 nsew signal output
rlabel metal2 s 23110 0 23166 800 6 wbs_dat_o[11]
port 574 nsew signal output
rlabel metal2 s 24582 0 24638 800 6 wbs_dat_o[12]
port 575 nsew signal output
rlabel metal2 s 26146 0 26202 800 6 wbs_dat_o[13]
port 576 nsew signal output
rlabel metal2 s 27618 0 27674 800 6 wbs_dat_o[14]
port 577 nsew signal output
rlabel metal2 s 29182 0 29238 800 6 wbs_dat_o[15]
port 578 nsew signal output
rlabel metal2 s 30746 0 30802 800 6 wbs_dat_o[16]
port 579 nsew signal output
rlabel metal2 s 32218 0 32274 800 6 wbs_dat_o[17]
port 580 nsew signal output
rlabel metal2 s 33782 0 33838 800 6 wbs_dat_o[18]
port 581 nsew signal output
rlabel metal2 s 35254 0 35310 800 6 wbs_dat_o[19]
port 582 nsew signal output
rlabel metal2 s 6274 0 6330 800 6 wbs_dat_o[1]
port 583 nsew signal output
rlabel metal2 s 36818 0 36874 800 6 wbs_dat_o[20]
port 584 nsew signal output
rlabel metal2 s 38382 0 38438 800 6 wbs_dat_o[21]
port 585 nsew signal output
rlabel metal2 s 39854 0 39910 800 6 wbs_dat_o[22]
port 586 nsew signal output
rlabel metal2 s 41418 0 41474 800 6 wbs_dat_o[23]
port 587 nsew signal output
rlabel metal2 s 42890 0 42946 800 6 wbs_dat_o[24]
port 588 nsew signal output
rlabel metal2 s 44454 0 44510 800 6 wbs_dat_o[25]
port 589 nsew signal output
rlabel metal2 s 46018 0 46074 800 6 wbs_dat_o[26]
port 590 nsew signal output
rlabel metal2 s 47490 0 47546 800 6 wbs_dat_o[27]
port 591 nsew signal output
rlabel metal2 s 49054 0 49110 800 6 wbs_dat_o[28]
port 592 nsew signal output
rlabel metal2 s 50526 0 50582 800 6 wbs_dat_o[29]
port 593 nsew signal output
rlabel metal2 s 8298 0 8354 800 6 wbs_dat_o[2]
port 594 nsew signal output
rlabel metal2 s 52090 0 52146 800 6 wbs_dat_o[30]
port 595 nsew signal output
rlabel metal2 s 53654 0 53710 800 6 wbs_dat_o[31]
port 596 nsew signal output
rlabel metal2 s 10322 0 10378 800 6 wbs_dat_o[3]
port 597 nsew signal output
rlabel metal2 s 12346 0 12402 800 6 wbs_dat_o[4]
port 598 nsew signal output
rlabel metal2 s 13910 0 13966 800 6 wbs_dat_o[5]
port 599 nsew signal output
rlabel metal2 s 15474 0 15530 800 6 wbs_dat_o[6]
port 600 nsew signal output
rlabel metal2 s 16946 0 17002 800 6 wbs_dat_o[7]
port 601 nsew signal output
rlabel metal2 s 18510 0 18566 800 6 wbs_dat_o[8]
port 602 nsew signal output
rlabel metal2 s 19982 0 20038 800 6 wbs_dat_o[9]
port 603 nsew signal output
rlabel metal2 s 4710 0 4766 800 6 wbs_sel_i[0]
port 604 nsew signal input
rlabel metal2 s 6734 0 6790 800 6 wbs_sel_i[1]
port 605 nsew signal input
rlabel metal2 s 8850 0 8906 800 6 wbs_sel_i[2]
port 606 nsew signal input
rlabel metal2 s 10874 0 10930 800 6 wbs_sel_i[3]
port 607 nsew signal input
rlabel metal2 s 2226 0 2282 800 6 wbs_stb_i
port 608 nsew signal input
rlabel metal2 s 2686 0 2742 800 6 wbs_we_i
port 609 nsew signal input
<< properties >>
string FIXED_BBOX 0 0 250000 250000
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 47646116
string GDS_FILE /home/fatihgulakar/638_proje/shooting_game_verilog/openlane/user_proj_example/runs/user_proj_example/results/finishing/user_proj_example.magic.gds
string GDS_START 1590158
<< end >>

