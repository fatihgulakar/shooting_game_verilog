module obj_heart  (
    input [3:0] x,
    input [3:0] y,
    input       en,
    output      data
);
    reg rom [0:14][0:14];
	
	initial begin
 rom[0][0] = 1'b0;	 rom[1][0] = 1'b0;	 rom[2][0] = 1'b0;	 rom[3][0] = 1'b0;	 rom[4][0] = 1'b0;	 rom[5][0] = 1'b0;	 rom[6][0] = 1'b0;	 rom[7][0] = 1'b0;	 rom[8][0] = 1'b0;	 rom[9][0] = 1'b0;	 rom[10][0] = 1'b0;	 rom[11][0] = 1'b0;	 rom[12][0] = 1'b0;	 rom[13][0] = 1'b0;	 rom[14][0] = 1'b0;
 rom[0][1] = 1'b0;	 rom[1][1] = 1'b0;	 rom[2][1] = 1'b0;	 rom[3][1] = 1'b0;	 rom[4][1] = 1'b0;	 rom[5][1] = 1'b0;	 rom[6][1] = 1'b0;	 rom[7][1] = 1'b0;	 rom[8][1] = 1'b0;	 rom[9][1] = 1'b0;	 rom[10][1] = 1'b0;	 rom[11][1] = 1'b0;	 rom[12][1] = 1'b0;	 rom[13][1] = 1'b0;	 rom[14][1] = 1'b0;
 rom[0][2] = 1'b0;	 rom[1][2] = 1'b0;	 rom[2][2] = 1'b0;	 rom[3][2] = 1'b1;	 rom[4][2] = 1'b1;	 rom[5][2] = 1'b1;	 rom[6][2] = 1'b0;	 rom[7][2] = 1'b0;	 rom[8][2] = 1'b0;	 rom[9][2] = 1'b1;	 rom[10][2] = 1'b1;	 rom[11][2] = 1'b1;	 rom[12][2] = 1'b0;	 rom[13][2] = 1'b0;	 rom[14][2] = 1'b0;
 rom[0][3] = 1'b0;	 rom[1][3] = 1'b0;	 rom[2][3] = 1'b1;	 rom[3][3] = 1'b0;	 rom[4][3] = 1'b0;	 rom[5][3] = 1'b1;	 rom[6][3] = 1'b1;	 rom[7][3] = 1'b0;	 rom[8][3] = 1'b1;	 rom[9][3] = 1'b1;	 rom[10][3] = 1'b1;	 rom[11][3] = 1'b1;	 rom[12][3] = 1'b1;	 rom[13][3] = 1'b0;	 rom[14][3] = 1'b0;
 rom[0][4] = 1'b0;	 rom[1][4] = 1'b1;	 rom[2][4] = 1'b0;	 rom[3][4] = 1'b0;	 rom[4][4] = 1'b1;	 rom[5][4] = 1'b1;	 rom[6][4] = 1'b1;	 rom[7][4] = 1'b1;	 rom[8][4] = 1'b1;	 rom[9][4] = 1'b1;	 rom[10][4] = 1'b1;	 rom[11][4] = 1'b1;	 rom[12][4] = 1'b1;	 rom[13][4] = 1'b1;	 rom[14][4] = 1'b0;
 rom[0][5] = 1'b0;	 rom[1][5] = 1'b1;	 rom[2][5] = 1'b1;	 rom[3][5] = 1'b1;	 rom[4][5] = 1'b1;	 rom[5][5] = 1'b1;	 rom[6][5] = 1'b1;	 rom[7][5] = 1'b1;	 rom[8][5] = 1'b1;	 rom[9][5] = 1'b1;	 rom[10][5] = 1'b1;	 rom[11][5] = 1'b1;	 rom[12][5] = 1'b1;	 rom[13][5] = 1'b1;	 rom[14][5] = 1'b0;
 rom[0][6] = 1'b0;	 rom[1][6] = 1'b1;	 rom[2][6] = 1'b1;	 rom[3][6] = 1'b1;	 rom[4][6] = 1'b1;	 rom[5][6] = 1'b1;	 rom[6][6] = 1'b1;	 rom[7][6] = 1'b1;	 rom[8][6] = 1'b1;	 rom[9][6] = 1'b1;	 rom[10][6] = 1'b1;	 rom[11][6] = 1'b1;	 rom[12][6] = 1'b1;	 rom[13][6] = 1'b1;	 rom[14][6] = 1'b0;
 rom[0][7] = 1'b0;	 rom[1][7] = 1'b0;	 rom[2][7] = 1'b1;	 rom[3][7] = 1'b1;	 rom[4][7] = 1'b1;	 rom[5][7] = 1'b1;	 rom[6][7] = 1'b1;	 rom[7][7] = 1'b1;	 rom[8][7] = 1'b1;	 rom[9][7] = 1'b1;	 rom[10][7] = 1'b1;	 rom[11][7] = 1'b1;	 rom[12][7] = 1'b1;	 rom[13][7] = 1'b0;	 rom[14][7] = 1'b0;
 rom[0][8] = 1'b0;	 rom[1][8] = 1'b0;	 rom[2][8] = 1'b0;	 rom[3][8] = 1'b1;	 rom[4][8] = 1'b1;	 rom[5][8] = 1'b1;	 rom[6][8] = 1'b1;	 rom[7][8] = 1'b1;	 rom[8][8] = 1'b1;	 rom[9][8] = 1'b1;	 rom[10][8] = 1'b1;	 rom[11][8] = 1'b1;	 rom[12][8] = 1'b0;	 rom[13][8] = 1'b0;	 rom[14][8] = 1'b0;
 rom[0][9] = 1'b0;	 rom[1][9] = 1'b0;	 rom[2][9] = 1'b0;	 rom[3][9] = 1'b0;	 rom[4][9] = 1'b1;	 rom[5][9] = 1'b1;	 rom[6][9] = 1'b1;	 rom[7][9] = 1'b1;	 rom[8][9] = 1'b1;	 rom[9][9] = 1'b1;	 rom[10][9] = 1'b1;	 rom[11][9] = 1'b0;	 rom[12][9] = 1'b0;	 rom[13][9] = 1'b0;	 rom[14][9] = 1'b0;
 rom[0][10] = 1'b0;	 rom[1][10] = 1'b0;	 rom[2][10] = 1'b0;	 rom[3][10] = 1'b0;	 rom[4][10] = 1'b0;	 rom[5][10] = 1'b1;	 rom[6][10] = 1'b1;	 rom[7][10] = 1'b1;	 rom[8][10] = 1'b1;	 rom[9][10] = 1'b1;	 rom[10][10] = 1'b0;	 rom[11][10] = 1'b0;	 rom[12][10] = 1'b0;	 rom[13][10] = 1'b0;	 rom[14][10] = 1'b0;
 rom[0][11] = 1'b0;	 rom[1][11] = 1'b0;	 rom[2][11] = 1'b0;	 rom[3][11] = 1'b0;	 rom[4][11] = 1'b0;	 rom[5][11] = 1'b0;	 rom[6][11] = 1'b1;	 rom[7][11] = 1'b1;	 rom[8][11] = 1'b1;	 rom[9][11] = 1'b0;	 rom[10][11] = 1'b0;	 rom[11][11] = 1'b0;	 rom[12][11] = 1'b0;	 rom[13][11] = 1'b0;	 rom[14][11] = 1'b0;
 rom[0][12] = 1'b0;	 rom[1][12] = 1'b0;	 rom[2][12] = 1'b0;	 rom[3][12] = 1'b0;	 rom[4][12] = 1'b0;	 rom[5][12] = 1'b0;	 rom[6][12] = 1'b0;	 rom[7][12] = 1'b1;	 rom[8][12] = 1'b0;	 rom[9][12] = 1'b0;	 rom[10][12] = 1'b0;	 rom[11][12] = 1'b0;	 rom[12][12] = 1'b0;	 rom[13][12] = 1'b0;	 rom[14][12] = 1'b0;
 rom[0][13] = 1'b0;	 rom[1][13] = 1'b0;	 rom[2][13] = 1'b0;	 rom[3][13] = 1'b0;	 rom[4][13] = 1'b0;	 rom[5][13] = 1'b0;	 rom[6][13] = 1'b0;	 rom[7][13] = 1'b0;	 rom[8][13] = 1'b0;	 rom[9][13] = 1'b0;	 rom[10][13] = 1'b0;	 rom[11][13] = 1'b0;	 rom[12][13] = 1'b0;	 rom[13][13] = 1'b0;	 rom[14][13] = 1'b0;
 rom[0][14] = 1'b0;	 rom[1][14] = 1'b0;	 rom[2][14] = 1'b0;	 rom[3][14] = 1'b0;	 rom[4][14] = 1'b0;	 rom[5][14] = 1'b0;	 rom[6][14] = 1'b0;	 rom[7][14] = 1'b0;	 rom[8][14] = 1'b0;	 rom[9][14] = 1'b0;	 rom[10][14] = 1'b0;	 rom[11][14] = 1'b0;	 rom[12][14] = 1'b0;	 rom[13][14] = 1'b0;	 rom[14][14] = 1'b0;
 end

    assign data = en ? rom[x][y] : 1'b0;

    
endmodule