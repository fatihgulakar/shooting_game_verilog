magic
tech sky130A
magscale 1 2
timestamp 1655299706
<< obsli1 >>
rect 1104 2159 248860 247537
<< obsm1 >>
rect 198 2128 249122 247568
<< metal2 >>
rect 4434 249200 4490 250000
rect 13358 249200 13414 250000
rect 22282 249200 22338 250000
rect 31206 249200 31262 250000
rect 40130 249200 40186 250000
rect 49054 249200 49110 250000
rect 57978 249200 58034 250000
rect 66902 249200 66958 250000
rect 75826 249200 75882 250000
rect 84750 249200 84806 250000
rect 93674 249200 93730 250000
rect 102598 249200 102654 250000
rect 111522 249200 111578 250000
rect 120446 249200 120502 250000
rect 129370 249200 129426 250000
rect 138294 249200 138350 250000
rect 147218 249200 147274 250000
rect 156142 249200 156198 250000
rect 165066 249200 165122 250000
rect 173990 249200 174046 250000
rect 182914 249200 182970 250000
rect 191838 249200 191894 250000
rect 200762 249200 200818 250000
rect 209686 249200 209742 250000
rect 218610 249200 218666 250000
rect 227534 249200 227590 250000
rect 236458 249200 236514 250000
rect 245382 249200 245438 250000
rect 202 0 258 800
rect 662 0 718 800
rect 1214 0 1270 800
rect 1674 0 1730 800
rect 2226 0 2282 800
rect 2686 0 2742 800
rect 3238 0 3294 800
rect 3698 0 3754 800
rect 4250 0 4306 800
rect 4710 0 4766 800
rect 5262 0 5318 800
rect 5722 0 5778 800
rect 6274 0 6330 800
rect 6826 0 6882 800
rect 7286 0 7342 800
rect 7838 0 7894 800
rect 8298 0 8354 800
rect 8850 0 8906 800
rect 9310 0 9366 800
rect 9862 0 9918 800
rect 10322 0 10378 800
rect 10874 0 10930 800
rect 11334 0 11390 800
rect 11886 0 11942 800
rect 12438 0 12494 800
rect 12898 0 12954 800
rect 13450 0 13506 800
rect 13910 0 13966 800
rect 14462 0 14518 800
rect 14922 0 14978 800
rect 15474 0 15530 800
rect 15934 0 15990 800
rect 16486 0 16542 800
rect 16946 0 17002 800
rect 17498 0 17554 800
rect 18050 0 18106 800
rect 18510 0 18566 800
rect 19062 0 19118 800
rect 19522 0 19578 800
rect 20074 0 20130 800
rect 20534 0 20590 800
rect 21086 0 21142 800
rect 21546 0 21602 800
rect 22098 0 22154 800
rect 22558 0 22614 800
rect 23110 0 23166 800
rect 23662 0 23718 800
rect 24122 0 24178 800
rect 24674 0 24730 800
rect 25134 0 25190 800
rect 25686 0 25742 800
rect 26146 0 26202 800
rect 26698 0 26754 800
rect 27158 0 27214 800
rect 27710 0 27766 800
rect 28170 0 28226 800
rect 28722 0 28778 800
rect 29274 0 29330 800
rect 29734 0 29790 800
rect 30286 0 30342 800
rect 30746 0 30802 800
rect 31298 0 31354 800
rect 31758 0 31814 800
rect 32310 0 32366 800
rect 32770 0 32826 800
rect 33322 0 33378 800
rect 33782 0 33838 800
rect 34334 0 34390 800
rect 34886 0 34942 800
rect 35346 0 35402 800
rect 35898 0 35954 800
rect 36358 0 36414 800
rect 36910 0 36966 800
rect 37370 0 37426 800
rect 37922 0 37978 800
rect 38382 0 38438 800
rect 38934 0 38990 800
rect 39394 0 39450 800
rect 39946 0 40002 800
rect 40498 0 40554 800
rect 40958 0 41014 800
rect 41510 0 41566 800
rect 41970 0 42026 800
rect 42522 0 42578 800
rect 42982 0 43038 800
rect 43534 0 43590 800
rect 43994 0 44050 800
rect 44546 0 44602 800
rect 45006 0 45062 800
rect 45558 0 45614 800
rect 46110 0 46166 800
rect 46570 0 46626 800
rect 47122 0 47178 800
rect 47582 0 47638 800
rect 48134 0 48190 800
rect 48594 0 48650 800
rect 49146 0 49202 800
rect 49606 0 49662 800
rect 50158 0 50214 800
rect 50618 0 50674 800
rect 51170 0 51226 800
rect 51722 0 51778 800
rect 52182 0 52238 800
rect 52734 0 52790 800
rect 53194 0 53250 800
rect 53746 0 53802 800
rect 54206 0 54262 800
rect 54758 0 54814 800
rect 55218 0 55274 800
rect 55770 0 55826 800
rect 56230 0 56286 800
rect 56782 0 56838 800
rect 57334 0 57390 800
rect 57794 0 57850 800
rect 58346 0 58402 800
rect 58806 0 58862 800
rect 59358 0 59414 800
rect 59818 0 59874 800
rect 60370 0 60426 800
rect 60830 0 60886 800
rect 61382 0 61438 800
rect 61842 0 61898 800
rect 62394 0 62450 800
rect 62946 0 63002 800
rect 63406 0 63462 800
rect 63958 0 64014 800
rect 64418 0 64474 800
rect 64970 0 65026 800
rect 65430 0 65486 800
rect 65982 0 66038 800
rect 66442 0 66498 800
rect 66994 0 67050 800
rect 67454 0 67510 800
rect 68006 0 68062 800
rect 68558 0 68614 800
rect 69018 0 69074 800
rect 69570 0 69626 800
rect 70030 0 70086 800
rect 70582 0 70638 800
rect 71042 0 71098 800
rect 71594 0 71650 800
rect 72054 0 72110 800
rect 72606 0 72662 800
rect 73066 0 73122 800
rect 73618 0 73674 800
rect 74170 0 74226 800
rect 74630 0 74686 800
rect 75182 0 75238 800
rect 75642 0 75698 800
rect 76194 0 76250 800
rect 76654 0 76710 800
rect 77206 0 77262 800
rect 77666 0 77722 800
rect 78218 0 78274 800
rect 78678 0 78734 800
rect 79230 0 79286 800
rect 79782 0 79838 800
rect 80242 0 80298 800
rect 80794 0 80850 800
rect 81254 0 81310 800
rect 81806 0 81862 800
rect 82266 0 82322 800
rect 82818 0 82874 800
rect 83278 0 83334 800
rect 83830 0 83886 800
rect 84290 0 84346 800
rect 84842 0 84898 800
rect 85302 0 85358 800
rect 85854 0 85910 800
rect 86406 0 86462 800
rect 86866 0 86922 800
rect 87418 0 87474 800
rect 87878 0 87934 800
rect 88430 0 88486 800
rect 88890 0 88946 800
rect 89442 0 89498 800
rect 89902 0 89958 800
rect 90454 0 90510 800
rect 90914 0 90970 800
rect 91466 0 91522 800
rect 92018 0 92074 800
rect 92478 0 92534 800
rect 93030 0 93086 800
rect 93490 0 93546 800
rect 94042 0 94098 800
rect 94502 0 94558 800
rect 95054 0 95110 800
rect 95514 0 95570 800
rect 96066 0 96122 800
rect 96526 0 96582 800
rect 97078 0 97134 800
rect 97630 0 97686 800
rect 98090 0 98146 800
rect 98642 0 98698 800
rect 99102 0 99158 800
rect 99654 0 99710 800
rect 100114 0 100170 800
rect 100666 0 100722 800
rect 101126 0 101182 800
rect 101678 0 101734 800
rect 102138 0 102194 800
rect 102690 0 102746 800
rect 103242 0 103298 800
rect 103702 0 103758 800
rect 104254 0 104310 800
rect 104714 0 104770 800
rect 105266 0 105322 800
rect 105726 0 105782 800
rect 106278 0 106334 800
rect 106738 0 106794 800
rect 107290 0 107346 800
rect 107750 0 107806 800
rect 108302 0 108358 800
rect 108854 0 108910 800
rect 109314 0 109370 800
rect 109866 0 109922 800
rect 110326 0 110382 800
rect 110878 0 110934 800
rect 111338 0 111394 800
rect 111890 0 111946 800
rect 112350 0 112406 800
rect 112902 0 112958 800
rect 113362 0 113418 800
rect 113914 0 113970 800
rect 114466 0 114522 800
rect 114926 0 114982 800
rect 115478 0 115534 800
rect 115938 0 115994 800
rect 116490 0 116546 800
rect 116950 0 117006 800
rect 117502 0 117558 800
rect 117962 0 118018 800
rect 118514 0 118570 800
rect 118974 0 119030 800
rect 119526 0 119582 800
rect 120078 0 120134 800
rect 120538 0 120594 800
rect 121090 0 121146 800
rect 121550 0 121606 800
rect 122102 0 122158 800
rect 122562 0 122618 800
rect 123114 0 123170 800
rect 123574 0 123630 800
rect 124126 0 124182 800
rect 124586 0 124642 800
rect 125138 0 125194 800
rect 125690 0 125746 800
rect 126150 0 126206 800
rect 126702 0 126758 800
rect 127162 0 127218 800
rect 127714 0 127770 800
rect 128174 0 128230 800
rect 128726 0 128782 800
rect 129186 0 129242 800
rect 129738 0 129794 800
rect 130198 0 130254 800
rect 130750 0 130806 800
rect 131302 0 131358 800
rect 131762 0 131818 800
rect 132314 0 132370 800
rect 132774 0 132830 800
rect 133326 0 133382 800
rect 133786 0 133842 800
rect 134338 0 134394 800
rect 134798 0 134854 800
rect 135350 0 135406 800
rect 135810 0 135866 800
rect 136362 0 136418 800
rect 136914 0 136970 800
rect 137374 0 137430 800
rect 137926 0 137982 800
rect 138386 0 138442 800
rect 138938 0 138994 800
rect 139398 0 139454 800
rect 139950 0 140006 800
rect 140410 0 140466 800
rect 140962 0 141018 800
rect 141422 0 141478 800
rect 141974 0 142030 800
rect 142526 0 142582 800
rect 142986 0 143042 800
rect 143538 0 143594 800
rect 143998 0 144054 800
rect 144550 0 144606 800
rect 145010 0 145066 800
rect 145562 0 145618 800
rect 146022 0 146078 800
rect 146574 0 146630 800
rect 147034 0 147090 800
rect 147586 0 147642 800
rect 148138 0 148194 800
rect 148598 0 148654 800
rect 149150 0 149206 800
rect 149610 0 149666 800
rect 150162 0 150218 800
rect 150622 0 150678 800
rect 151174 0 151230 800
rect 151634 0 151690 800
rect 152186 0 152242 800
rect 152646 0 152702 800
rect 153198 0 153254 800
rect 153750 0 153806 800
rect 154210 0 154266 800
rect 154762 0 154818 800
rect 155222 0 155278 800
rect 155774 0 155830 800
rect 156234 0 156290 800
rect 156786 0 156842 800
rect 157246 0 157302 800
rect 157798 0 157854 800
rect 158258 0 158314 800
rect 158810 0 158866 800
rect 159362 0 159418 800
rect 159822 0 159878 800
rect 160374 0 160430 800
rect 160834 0 160890 800
rect 161386 0 161442 800
rect 161846 0 161902 800
rect 162398 0 162454 800
rect 162858 0 162914 800
rect 163410 0 163466 800
rect 163870 0 163926 800
rect 164422 0 164478 800
rect 164974 0 165030 800
rect 165434 0 165490 800
rect 165986 0 166042 800
rect 166446 0 166502 800
rect 166998 0 167054 800
rect 167458 0 167514 800
rect 168010 0 168066 800
rect 168470 0 168526 800
rect 169022 0 169078 800
rect 169482 0 169538 800
rect 170034 0 170090 800
rect 170494 0 170550 800
rect 171046 0 171102 800
rect 171598 0 171654 800
rect 172058 0 172114 800
rect 172610 0 172666 800
rect 173070 0 173126 800
rect 173622 0 173678 800
rect 174082 0 174138 800
rect 174634 0 174690 800
rect 175094 0 175150 800
rect 175646 0 175702 800
rect 176106 0 176162 800
rect 176658 0 176714 800
rect 177210 0 177266 800
rect 177670 0 177726 800
rect 178222 0 178278 800
rect 178682 0 178738 800
rect 179234 0 179290 800
rect 179694 0 179750 800
rect 180246 0 180302 800
rect 180706 0 180762 800
rect 181258 0 181314 800
rect 181718 0 181774 800
rect 182270 0 182326 800
rect 182822 0 182878 800
rect 183282 0 183338 800
rect 183834 0 183890 800
rect 184294 0 184350 800
rect 184846 0 184902 800
rect 185306 0 185362 800
rect 185858 0 185914 800
rect 186318 0 186374 800
rect 186870 0 186926 800
rect 187330 0 187386 800
rect 187882 0 187938 800
rect 188434 0 188490 800
rect 188894 0 188950 800
rect 189446 0 189502 800
rect 189906 0 189962 800
rect 190458 0 190514 800
rect 190918 0 190974 800
rect 191470 0 191526 800
rect 191930 0 191986 800
rect 192482 0 192538 800
rect 192942 0 192998 800
rect 193494 0 193550 800
rect 194046 0 194102 800
rect 194506 0 194562 800
rect 195058 0 195114 800
rect 195518 0 195574 800
rect 196070 0 196126 800
rect 196530 0 196586 800
rect 197082 0 197138 800
rect 197542 0 197598 800
rect 198094 0 198150 800
rect 198554 0 198610 800
rect 199106 0 199162 800
rect 199658 0 199714 800
rect 200118 0 200174 800
rect 200670 0 200726 800
rect 201130 0 201186 800
rect 201682 0 201738 800
rect 202142 0 202198 800
rect 202694 0 202750 800
rect 203154 0 203210 800
rect 203706 0 203762 800
rect 204166 0 204222 800
rect 204718 0 204774 800
rect 205270 0 205326 800
rect 205730 0 205786 800
rect 206282 0 206338 800
rect 206742 0 206798 800
rect 207294 0 207350 800
rect 207754 0 207810 800
rect 208306 0 208362 800
rect 208766 0 208822 800
rect 209318 0 209374 800
rect 209778 0 209834 800
rect 210330 0 210386 800
rect 210882 0 210938 800
rect 211342 0 211398 800
rect 211894 0 211950 800
rect 212354 0 212410 800
rect 212906 0 212962 800
rect 213366 0 213422 800
rect 213918 0 213974 800
rect 214378 0 214434 800
rect 214930 0 214986 800
rect 215390 0 215446 800
rect 215942 0 215998 800
rect 216494 0 216550 800
rect 216954 0 217010 800
rect 217506 0 217562 800
rect 217966 0 218022 800
rect 218518 0 218574 800
rect 218978 0 219034 800
rect 219530 0 219586 800
rect 219990 0 220046 800
rect 220542 0 220598 800
rect 221002 0 221058 800
rect 221554 0 221610 800
rect 222106 0 222162 800
rect 222566 0 222622 800
rect 223118 0 223174 800
rect 223578 0 223634 800
rect 224130 0 224186 800
rect 224590 0 224646 800
rect 225142 0 225198 800
rect 225602 0 225658 800
rect 226154 0 226210 800
rect 226614 0 226670 800
rect 227166 0 227222 800
rect 227718 0 227774 800
rect 228178 0 228234 800
rect 228730 0 228786 800
rect 229190 0 229246 800
rect 229742 0 229798 800
rect 230202 0 230258 800
rect 230754 0 230810 800
rect 231214 0 231270 800
rect 231766 0 231822 800
rect 232226 0 232282 800
rect 232778 0 232834 800
rect 233330 0 233386 800
rect 233790 0 233846 800
rect 234342 0 234398 800
rect 234802 0 234858 800
rect 235354 0 235410 800
rect 235814 0 235870 800
rect 236366 0 236422 800
rect 236826 0 236882 800
rect 237378 0 237434 800
rect 237838 0 237894 800
rect 238390 0 238446 800
rect 238942 0 238998 800
rect 239402 0 239458 800
rect 239954 0 240010 800
rect 240414 0 240470 800
rect 240966 0 241022 800
rect 241426 0 241482 800
rect 241978 0 242034 800
rect 242438 0 242494 800
rect 242990 0 243046 800
rect 243450 0 243506 800
rect 244002 0 244058 800
rect 244554 0 244610 800
rect 245014 0 245070 800
rect 245566 0 245622 800
rect 246026 0 246082 800
rect 246578 0 246634 800
rect 247038 0 247094 800
rect 247590 0 247646 800
rect 248050 0 248106 800
rect 248602 0 248658 800
rect 249062 0 249118 800
rect 249614 0 249670 800
<< obsm2 >>
rect 204 249144 4378 249234
rect 4546 249144 13302 249234
rect 13470 249144 22226 249234
rect 22394 249144 31150 249234
rect 31318 249144 40074 249234
rect 40242 249144 48998 249234
rect 49166 249144 57922 249234
rect 58090 249144 66846 249234
rect 67014 249144 75770 249234
rect 75938 249144 84694 249234
rect 84862 249144 93618 249234
rect 93786 249144 102542 249234
rect 102710 249144 111466 249234
rect 111634 249144 120390 249234
rect 120558 249144 129314 249234
rect 129482 249144 138238 249234
rect 138406 249144 147162 249234
rect 147330 249144 156086 249234
rect 156254 249144 165010 249234
rect 165178 249144 173934 249234
rect 174102 249144 182858 249234
rect 183026 249144 191782 249234
rect 191950 249144 200706 249234
rect 200874 249144 209630 249234
rect 209798 249144 218554 249234
rect 218722 249144 227478 249234
rect 227646 249144 236402 249234
rect 236570 249144 245326 249234
rect 245494 249144 249116 249234
rect 204 856 249116 249144
rect 314 800 606 856
rect 774 800 1158 856
rect 1326 800 1618 856
rect 1786 800 2170 856
rect 2338 800 2630 856
rect 2798 800 3182 856
rect 3350 800 3642 856
rect 3810 800 4194 856
rect 4362 800 4654 856
rect 4822 800 5206 856
rect 5374 800 5666 856
rect 5834 800 6218 856
rect 6386 800 6770 856
rect 6938 800 7230 856
rect 7398 800 7782 856
rect 7950 800 8242 856
rect 8410 800 8794 856
rect 8962 800 9254 856
rect 9422 800 9806 856
rect 9974 800 10266 856
rect 10434 800 10818 856
rect 10986 800 11278 856
rect 11446 800 11830 856
rect 11998 800 12382 856
rect 12550 800 12842 856
rect 13010 800 13394 856
rect 13562 800 13854 856
rect 14022 800 14406 856
rect 14574 800 14866 856
rect 15034 800 15418 856
rect 15586 800 15878 856
rect 16046 800 16430 856
rect 16598 800 16890 856
rect 17058 800 17442 856
rect 17610 800 17994 856
rect 18162 800 18454 856
rect 18622 800 19006 856
rect 19174 800 19466 856
rect 19634 800 20018 856
rect 20186 800 20478 856
rect 20646 800 21030 856
rect 21198 800 21490 856
rect 21658 800 22042 856
rect 22210 800 22502 856
rect 22670 800 23054 856
rect 23222 800 23606 856
rect 23774 800 24066 856
rect 24234 800 24618 856
rect 24786 800 25078 856
rect 25246 800 25630 856
rect 25798 800 26090 856
rect 26258 800 26642 856
rect 26810 800 27102 856
rect 27270 800 27654 856
rect 27822 800 28114 856
rect 28282 800 28666 856
rect 28834 800 29218 856
rect 29386 800 29678 856
rect 29846 800 30230 856
rect 30398 800 30690 856
rect 30858 800 31242 856
rect 31410 800 31702 856
rect 31870 800 32254 856
rect 32422 800 32714 856
rect 32882 800 33266 856
rect 33434 800 33726 856
rect 33894 800 34278 856
rect 34446 800 34830 856
rect 34998 800 35290 856
rect 35458 800 35842 856
rect 36010 800 36302 856
rect 36470 800 36854 856
rect 37022 800 37314 856
rect 37482 800 37866 856
rect 38034 800 38326 856
rect 38494 800 38878 856
rect 39046 800 39338 856
rect 39506 800 39890 856
rect 40058 800 40442 856
rect 40610 800 40902 856
rect 41070 800 41454 856
rect 41622 800 41914 856
rect 42082 800 42466 856
rect 42634 800 42926 856
rect 43094 800 43478 856
rect 43646 800 43938 856
rect 44106 800 44490 856
rect 44658 800 44950 856
rect 45118 800 45502 856
rect 45670 800 46054 856
rect 46222 800 46514 856
rect 46682 800 47066 856
rect 47234 800 47526 856
rect 47694 800 48078 856
rect 48246 800 48538 856
rect 48706 800 49090 856
rect 49258 800 49550 856
rect 49718 800 50102 856
rect 50270 800 50562 856
rect 50730 800 51114 856
rect 51282 800 51666 856
rect 51834 800 52126 856
rect 52294 800 52678 856
rect 52846 800 53138 856
rect 53306 800 53690 856
rect 53858 800 54150 856
rect 54318 800 54702 856
rect 54870 800 55162 856
rect 55330 800 55714 856
rect 55882 800 56174 856
rect 56342 800 56726 856
rect 56894 800 57278 856
rect 57446 800 57738 856
rect 57906 800 58290 856
rect 58458 800 58750 856
rect 58918 800 59302 856
rect 59470 800 59762 856
rect 59930 800 60314 856
rect 60482 800 60774 856
rect 60942 800 61326 856
rect 61494 800 61786 856
rect 61954 800 62338 856
rect 62506 800 62890 856
rect 63058 800 63350 856
rect 63518 800 63902 856
rect 64070 800 64362 856
rect 64530 800 64914 856
rect 65082 800 65374 856
rect 65542 800 65926 856
rect 66094 800 66386 856
rect 66554 800 66938 856
rect 67106 800 67398 856
rect 67566 800 67950 856
rect 68118 800 68502 856
rect 68670 800 68962 856
rect 69130 800 69514 856
rect 69682 800 69974 856
rect 70142 800 70526 856
rect 70694 800 70986 856
rect 71154 800 71538 856
rect 71706 800 71998 856
rect 72166 800 72550 856
rect 72718 800 73010 856
rect 73178 800 73562 856
rect 73730 800 74114 856
rect 74282 800 74574 856
rect 74742 800 75126 856
rect 75294 800 75586 856
rect 75754 800 76138 856
rect 76306 800 76598 856
rect 76766 800 77150 856
rect 77318 800 77610 856
rect 77778 800 78162 856
rect 78330 800 78622 856
rect 78790 800 79174 856
rect 79342 800 79726 856
rect 79894 800 80186 856
rect 80354 800 80738 856
rect 80906 800 81198 856
rect 81366 800 81750 856
rect 81918 800 82210 856
rect 82378 800 82762 856
rect 82930 800 83222 856
rect 83390 800 83774 856
rect 83942 800 84234 856
rect 84402 800 84786 856
rect 84954 800 85246 856
rect 85414 800 85798 856
rect 85966 800 86350 856
rect 86518 800 86810 856
rect 86978 800 87362 856
rect 87530 800 87822 856
rect 87990 800 88374 856
rect 88542 800 88834 856
rect 89002 800 89386 856
rect 89554 800 89846 856
rect 90014 800 90398 856
rect 90566 800 90858 856
rect 91026 800 91410 856
rect 91578 800 91962 856
rect 92130 800 92422 856
rect 92590 800 92974 856
rect 93142 800 93434 856
rect 93602 800 93986 856
rect 94154 800 94446 856
rect 94614 800 94998 856
rect 95166 800 95458 856
rect 95626 800 96010 856
rect 96178 800 96470 856
rect 96638 800 97022 856
rect 97190 800 97574 856
rect 97742 800 98034 856
rect 98202 800 98586 856
rect 98754 800 99046 856
rect 99214 800 99598 856
rect 99766 800 100058 856
rect 100226 800 100610 856
rect 100778 800 101070 856
rect 101238 800 101622 856
rect 101790 800 102082 856
rect 102250 800 102634 856
rect 102802 800 103186 856
rect 103354 800 103646 856
rect 103814 800 104198 856
rect 104366 800 104658 856
rect 104826 800 105210 856
rect 105378 800 105670 856
rect 105838 800 106222 856
rect 106390 800 106682 856
rect 106850 800 107234 856
rect 107402 800 107694 856
rect 107862 800 108246 856
rect 108414 800 108798 856
rect 108966 800 109258 856
rect 109426 800 109810 856
rect 109978 800 110270 856
rect 110438 800 110822 856
rect 110990 800 111282 856
rect 111450 800 111834 856
rect 112002 800 112294 856
rect 112462 800 112846 856
rect 113014 800 113306 856
rect 113474 800 113858 856
rect 114026 800 114410 856
rect 114578 800 114870 856
rect 115038 800 115422 856
rect 115590 800 115882 856
rect 116050 800 116434 856
rect 116602 800 116894 856
rect 117062 800 117446 856
rect 117614 800 117906 856
rect 118074 800 118458 856
rect 118626 800 118918 856
rect 119086 800 119470 856
rect 119638 800 120022 856
rect 120190 800 120482 856
rect 120650 800 121034 856
rect 121202 800 121494 856
rect 121662 800 122046 856
rect 122214 800 122506 856
rect 122674 800 123058 856
rect 123226 800 123518 856
rect 123686 800 124070 856
rect 124238 800 124530 856
rect 124698 800 125082 856
rect 125250 800 125634 856
rect 125802 800 126094 856
rect 126262 800 126646 856
rect 126814 800 127106 856
rect 127274 800 127658 856
rect 127826 800 128118 856
rect 128286 800 128670 856
rect 128838 800 129130 856
rect 129298 800 129682 856
rect 129850 800 130142 856
rect 130310 800 130694 856
rect 130862 800 131246 856
rect 131414 800 131706 856
rect 131874 800 132258 856
rect 132426 800 132718 856
rect 132886 800 133270 856
rect 133438 800 133730 856
rect 133898 800 134282 856
rect 134450 800 134742 856
rect 134910 800 135294 856
rect 135462 800 135754 856
rect 135922 800 136306 856
rect 136474 800 136858 856
rect 137026 800 137318 856
rect 137486 800 137870 856
rect 138038 800 138330 856
rect 138498 800 138882 856
rect 139050 800 139342 856
rect 139510 800 139894 856
rect 140062 800 140354 856
rect 140522 800 140906 856
rect 141074 800 141366 856
rect 141534 800 141918 856
rect 142086 800 142470 856
rect 142638 800 142930 856
rect 143098 800 143482 856
rect 143650 800 143942 856
rect 144110 800 144494 856
rect 144662 800 144954 856
rect 145122 800 145506 856
rect 145674 800 145966 856
rect 146134 800 146518 856
rect 146686 800 146978 856
rect 147146 800 147530 856
rect 147698 800 148082 856
rect 148250 800 148542 856
rect 148710 800 149094 856
rect 149262 800 149554 856
rect 149722 800 150106 856
rect 150274 800 150566 856
rect 150734 800 151118 856
rect 151286 800 151578 856
rect 151746 800 152130 856
rect 152298 800 152590 856
rect 152758 800 153142 856
rect 153310 800 153694 856
rect 153862 800 154154 856
rect 154322 800 154706 856
rect 154874 800 155166 856
rect 155334 800 155718 856
rect 155886 800 156178 856
rect 156346 800 156730 856
rect 156898 800 157190 856
rect 157358 800 157742 856
rect 157910 800 158202 856
rect 158370 800 158754 856
rect 158922 800 159306 856
rect 159474 800 159766 856
rect 159934 800 160318 856
rect 160486 800 160778 856
rect 160946 800 161330 856
rect 161498 800 161790 856
rect 161958 800 162342 856
rect 162510 800 162802 856
rect 162970 800 163354 856
rect 163522 800 163814 856
rect 163982 800 164366 856
rect 164534 800 164918 856
rect 165086 800 165378 856
rect 165546 800 165930 856
rect 166098 800 166390 856
rect 166558 800 166942 856
rect 167110 800 167402 856
rect 167570 800 167954 856
rect 168122 800 168414 856
rect 168582 800 168966 856
rect 169134 800 169426 856
rect 169594 800 169978 856
rect 170146 800 170438 856
rect 170606 800 170990 856
rect 171158 800 171542 856
rect 171710 800 172002 856
rect 172170 800 172554 856
rect 172722 800 173014 856
rect 173182 800 173566 856
rect 173734 800 174026 856
rect 174194 800 174578 856
rect 174746 800 175038 856
rect 175206 800 175590 856
rect 175758 800 176050 856
rect 176218 800 176602 856
rect 176770 800 177154 856
rect 177322 800 177614 856
rect 177782 800 178166 856
rect 178334 800 178626 856
rect 178794 800 179178 856
rect 179346 800 179638 856
rect 179806 800 180190 856
rect 180358 800 180650 856
rect 180818 800 181202 856
rect 181370 800 181662 856
rect 181830 800 182214 856
rect 182382 800 182766 856
rect 182934 800 183226 856
rect 183394 800 183778 856
rect 183946 800 184238 856
rect 184406 800 184790 856
rect 184958 800 185250 856
rect 185418 800 185802 856
rect 185970 800 186262 856
rect 186430 800 186814 856
rect 186982 800 187274 856
rect 187442 800 187826 856
rect 187994 800 188378 856
rect 188546 800 188838 856
rect 189006 800 189390 856
rect 189558 800 189850 856
rect 190018 800 190402 856
rect 190570 800 190862 856
rect 191030 800 191414 856
rect 191582 800 191874 856
rect 192042 800 192426 856
rect 192594 800 192886 856
rect 193054 800 193438 856
rect 193606 800 193990 856
rect 194158 800 194450 856
rect 194618 800 195002 856
rect 195170 800 195462 856
rect 195630 800 196014 856
rect 196182 800 196474 856
rect 196642 800 197026 856
rect 197194 800 197486 856
rect 197654 800 198038 856
rect 198206 800 198498 856
rect 198666 800 199050 856
rect 199218 800 199602 856
rect 199770 800 200062 856
rect 200230 800 200614 856
rect 200782 800 201074 856
rect 201242 800 201626 856
rect 201794 800 202086 856
rect 202254 800 202638 856
rect 202806 800 203098 856
rect 203266 800 203650 856
rect 203818 800 204110 856
rect 204278 800 204662 856
rect 204830 800 205214 856
rect 205382 800 205674 856
rect 205842 800 206226 856
rect 206394 800 206686 856
rect 206854 800 207238 856
rect 207406 800 207698 856
rect 207866 800 208250 856
rect 208418 800 208710 856
rect 208878 800 209262 856
rect 209430 800 209722 856
rect 209890 800 210274 856
rect 210442 800 210826 856
rect 210994 800 211286 856
rect 211454 800 211838 856
rect 212006 800 212298 856
rect 212466 800 212850 856
rect 213018 800 213310 856
rect 213478 800 213862 856
rect 214030 800 214322 856
rect 214490 800 214874 856
rect 215042 800 215334 856
rect 215502 800 215886 856
rect 216054 800 216438 856
rect 216606 800 216898 856
rect 217066 800 217450 856
rect 217618 800 217910 856
rect 218078 800 218462 856
rect 218630 800 218922 856
rect 219090 800 219474 856
rect 219642 800 219934 856
rect 220102 800 220486 856
rect 220654 800 220946 856
rect 221114 800 221498 856
rect 221666 800 222050 856
rect 222218 800 222510 856
rect 222678 800 223062 856
rect 223230 800 223522 856
rect 223690 800 224074 856
rect 224242 800 224534 856
rect 224702 800 225086 856
rect 225254 800 225546 856
rect 225714 800 226098 856
rect 226266 800 226558 856
rect 226726 800 227110 856
rect 227278 800 227662 856
rect 227830 800 228122 856
rect 228290 800 228674 856
rect 228842 800 229134 856
rect 229302 800 229686 856
rect 229854 800 230146 856
rect 230314 800 230698 856
rect 230866 800 231158 856
rect 231326 800 231710 856
rect 231878 800 232170 856
rect 232338 800 232722 856
rect 232890 800 233274 856
rect 233442 800 233734 856
rect 233902 800 234286 856
rect 234454 800 234746 856
rect 234914 800 235298 856
rect 235466 800 235758 856
rect 235926 800 236310 856
rect 236478 800 236770 856
rect 236938 800 237322 856
rect 237490 800 237782 856
rect 237950 800 238334 856
rect 238502 800 238886 856
rect 239054 800 239346 856
rect 239514 800 239898 856
rect 240066 800 240358 856
rect 240526 800 240910 856
rect 241078 800 241370 856
rect 241538 800 241922 856
rect 242090 800 242382 856
rect 242550 800 242934 856
rect 243102 800 243394 856
rect 243562 800 243946 856
rect 244114 800 244498 856
rect 244666 800 244958 856
rect 245126 800 245510 856
rect 245678 800 245970 856
rect 246138 800 246522 856
rect 246690 800 246982 856
rect 247150 800 247534 856
rect 247702 800 247994 856
rect 248162 800 248546 856
rect 248714 800 249006 856
<< metal3 >>
rect 0 246984 800 247104
rect 249200 247120 250000 247240
rect 249200 241544 250000 241664
rect 0 241272 800 241392
rect 249200 235968 250000 236088
rect 0 235560 800 235680
rect 249200 230392 250000 230512
rect 0 229848 800 229968
rect 249200 224816 250000 224936
rect 0 224272 800 224392
rect 249200 219240 250000 219360
rect 0 218560 800 218680
rect 249200 213800 250000 213920
rect 0 212848 800 212968
rect 249200 208224 250000 208344
rect 0 207136 800 207256
rect 249200 202648 250000 202768
rect 0 201560 800 201680
rect 249200 197072 250000 197192
rect 0 195848 800 195968
rect 249200 191496 250000 191616
rect 0 190136 800 190256
rect 249200 185920 250000 186040
rect 0 184424 800 184544
rect 249200 180480 250000 180600
rect 0 178712 800 178832
rect 249200 174904 250000 175024
rect 0 173136 800 173256
rect 249200 169328 250000 169448
rect 0 167424 800 167544
rect 249200 163752 250000 163872
rect 0 161712 800 161832
rect 249200 158176 250000 158296
rect 0 156000 800 156120
rect 249200 152600 250000 152720
rect 0 150424 800 150544
rect 249200 147024 250000 147144
rect 0 144712 800 144832
rect 249200 141584 250000 141704
rect 0 139000 800 139120
rect 249200 136008 250000 136128
rect 0 133288 800 133408
rect 249200 130432 250000 130552
rect 0 127712 800 127832
rect 249200 124856 250000 124976
rect 0 122000 800 122120
rect 249200 119280 250000 119400
rect 0 116288 800 116408
rect 249200 113704 250000 113824
rect 0 110576 800 110696
rect 249200 108264 250000 108384
rect 0 104864 800 104984
rect 249200 102688 250000 102808
rect 0 99288 800 99408
rect 249200 97112 250000 97232
rect 0 93576 800 93696
rect 249200 91536 250000 91656
rect 0 87864 800 87984
rect 249200 85960 250000 86080
rect 0 82152 800 82272
rect 249200 80384 250000 80504
rect 0 76576 800 76696
rect 249200 74808 250000 74928
rect 0 70864 800 70984
rect 249200 69368 250000 69488
rect 0 65152 800 65272
rect 249200 63792 250000 63912
rect 0 59440 800 59560
rect 249200 58216 250000 58336
rect 0 53728 800 53848
rect 249200 52640 250000 52760
rect 0 48152 800 48272
rect 249200 47064 250000 47184
rect 0 42440 800 42560
rect 249200 41488 250000 41608
rect 0 36728 800 36848
rect 249200 36048 250000 36168
rect 0 31016 800 31136
rect 249200 30472 250000 30592
rect 0 25440 800 25560
rect 249200 24896 250000 25016
rect 0 19728 800 19848
rect 249200 19320 250000 19440
rect 0 14016 800 14136
rect 249200 13744 250000 13864
rect 0 8304 800 8424
rect 249200 8168 250000 8288
rect 0 2728 800 2848
rect 249200 2728 250000 2848
<< obsm3 >>
rect 800 247320 249200 247553
rect 800 247184 249120 247320
rect 880 247040 249120 247184
rect 880 246904 249200 247040
rect 800 241744 249200 246904
rect 800 241472 249120 241744
rect 880 241464 249120 241472
rect 880 241192 249200 241464
rect 800 236168 249200 241192
rect 800 235888 249120 236168
rect 800 235760 249200 235888
rect 880 235480 249200 235760
rect 800 230592 249200 235480
rect 800 230312 249120 230592
rect 800 230048 249200 230312
rect 880 229768 249200 230048
rect 800 225016 249200 229768
rect 800 224736 249120 225016
rect 800 224472 249200 224736
rect 880 224192 249200 224472
rect 800 219440 249200 224192
rect 800 219160 249120 219440
rect 800 218760 249200 219160
rect 880 218480 249200 218760
rect 800 214000 249200 218480
rect 800 213720 249120 214000
rect 800 213048 249200 213720
rect 880 212768 249200 213048
rect 800 208424 249200 212768
rect 800 208144 249120 208424
rect 800 207336 249200 208144
rect 880 207056 249200 207336
rect 800 202848 249200 207056
rect 800 202568 249120 202848
rect 800 201760 249200 202568
rect 880 201480 249200 201760
rect 800 197272 249200 201480
rect 800 196992 249120 197272
rect 800 196048 249200 196992
rect 880 195768 249200 196048
rect 800 191696 249200 195768
rect 800 191416 249120 191696
rect 800 190336 249200 191416
rect 880 190056 249200 190336
rect 800 186120 249200 190056
rect 800 185840 249120 186120
rect 800 184624 249200 185840
rect 880 184344 249200 184624
rect 800 180680 249200 184344
rect 800 180400 249120 180680
rect 800 178912 249200 180400
rect 880 178632 249200 178912
rect 800 175104 249200 178632
rect 800 174824 249120 175104
rect 800 173336 249200 174824
rect 880 173056 249200 173336
rect 800 169528 249200 173056
rect 800 169248 249120 169528
rect 800 167624 249200 169248
rect 880 167344 249200 167624
rect 800 163952 249200 167344
rect 800 163672 249120 163952
rect 800 161912 249200 163672
rect 880 161632 249200 161912
rect 800 158376 249200 161632
rect 800 158096 249120 158376
rect 800 156200 249200 158096
rect 880 155920 249200 156200
rect 800 152800 249200 155920
rect 800 152520 249120 152800
rect 800 150624 249200 152520
rect 880 150344 249200 150624
rect 800 147224 249200 150344
rect 800 146944 249120 147224
rect 800 144912 249200 146944
rect 880 144632 249200 144912
rect 800 141784 249200 144632
rect 800 141504 249120 141784
rect 800 139200 249200 141504
rect 880 138920 249200 139200
rect 800 136208 249200 138920
rect 800 135928 249120 136208
rect 800 133488 249200 135928
rect 880 133208 249200 133488
rect 800 130632 249200 133208
rect 800 130352 249120 130632
rect 800 127912 249200 130352
rect 880 127632 249200 127912
rect 800 125056 249200 127632
rect 800 124776 249120 125056
rect 800 122200 249200 124776
rect 880 121920 249200 122200
rect 800 119480 249200 121920
rect 800 119200 249120 119480
rect 800 116488 249200 119200
rect 880 116208 249200 116488
rect 800 113904 249200 116208
rect 800 113624 249120 113904
rect 800 110776 249200 113624
rect 880 110496 249200 110776
rect 800 108464 249200 110496
rect 800 108184 249120 108464
rect 800 105064 249200 108184
rect 880 104784 249200 105064
rect 800 102888 249200 104784
rect 800 102608 249120 102888
rect 800 99488 249200 102608
rect 880 99208 249200 99488
rect 800 97312 249200 99208
rect 800 97032 249120 97312
rect 800 93776 249200 97032
rect 880 93496 249200 93776
rect 800 91736 249200 93496
rect 800 91456 249120 91736
rect 800 88064 249200 91456
rect 880 87784 249200 88064
rect 800 86160 249200 87784
rect 800 85880 249120 86160
rect 800 82352 249200 85880
rect 880 82072 249200 82352
rect 800 80584 249200 82072
rect 800 80304 249120 80584
rect 800 76776 249200 80304
rect 880 76496 249200 76776
rect 800 75008 249200 76496
rect 800 74728 249120 75008
rect 800 71064 249200 74728
rect 880 70784 249200 71064
rect 800 69568 249200 70784
rect 800 69288 249120 69568
rect 800 65352 249200 69288
rect 880 65072 249200 65352
rect 800 63992 249200 65072
rect 800 63712 249120 63992
rect 800 59640 249200 63712
rect 880 59360 249200 59640
rect 800 58416 249200 59360
rect 800 58136 249120 58416
rect 800 53928 249200 58136
rect 880 53648 249200 53928
rect 800 52840 249200 53648
rect 800 52560 249120 52840
rect 800 48352 249200 52560
rect 880 48072 249200 48352
rect 800 47264 249200 48072
rect 800 46984 249120 47264
rect 800 42640 249200 46984
rect 880 42360 249200 42640
rect 800 41688 249200 42360
rect 800 41408 249120 41688
rect 800 36928 249200 41408
rect 880 36648 249200 36928
rect 800 36248 249200 36648
rect 800 35968 249120 36248
rect 800 31216 249200 35968
rect 880 30936 249200 31216
rect 800 30672 249200 30936
rect 800 30392 249120 30672
rect 800 25640 249200 30392
rect 880 25360 249200 25640
rect 800 25096 249200 25360
rect 800 24816 249120 25096
rect 800 19928 249200 24816
rect 880 19648 249200 19928
rect 800 19520 249200 19648
rect 800 19240 249120 19520
rect 800 14216 249200 19240
rect 880 13944 249200 14216
rect 880 13936 249120 13944
rect 800 13664 249120 13936
rect 800 8504 249200 13664
rect 880 8368 249200 8504
rect 880 8224 249120 8368
rect 800 8088 249120 8224
rect 800 2928 249200 8088
rect 880 2648 249120 2928
rect 800 2143 249200 2648
<< metal4 >>
rect 4208 2128 4528 247568
rect 19568 2128 19888 247568
rect 34928 2128 35248 247568
rect 50288 2128 50608 247568
rect 65648 2128 65968 247568
rect 81008 2128 81328 247568
rect 96368 2128 96688 247568
rect 111728 2128 112048 247568
rect 127088 2128 127408 247568
rect 142448 2128 142768 247568
rect 157808 2128 158128 247568
rect 173168 2128 173488 247568
rect 188528 2128 188848 247568
rect 203888 2128 204208 247568
rect 219248 2128 219568 247568
rect 234608 2128 234928 247568
<< obsm4 >>
rect 64275 2619 65568 162213
rect 66048 2619 80928 162213
rect 81408 2619 96288 162213
rect 96768 2619 111648 162213
rect 112128 2619 127008 162213
rect 127488 2619 142368 162213
rect 142848 2619 157728 162213
rect 158208 2619 173088 162213
rect 173568 2619 188448 162213
rect 188928 2619 202709 162213
<< labels >>
rlabel metal3 s 249200 2728 250000 2848 6 io_in[0]
port 1 nsew signal input
rlabel metal3 s 249200 169328 250000 169448 6 io_in[10]
port 2 nsew signal input
rlabel metal3 s 249200 185920 250000 186040 6 io_in[11]
port 3 nsew signal input
rlabel metal3 s 249200 202648 250000 202768 6 io_in[12]
port 4 nsew signal input
rlabel metal3 s 249200 219240 250000 219360 6 io_in[13]
port 5 nsew signal input
rlabel metal3 s 249200 235968 250000 236088 6 io_in[14]
port 6 nsew signal input
rlabel metal2 s 245382 249200 245438 250000 6 io_in[15]
port 7 nsew signal input
rlabel metal2 s 218610 249200 218666 250000 6 io_in[16]
port 8 nsew signal input
rlabel metal2 s 191838 249200 191894 250000 6 io_in[17]
port 9 nsew signal input
rlabel metal2 s 165066 249200 165122 250000 6 io_in[18]
port 10 nsew signal input
rlabel metal2 s 138294 249200 138350 250000 6 io_in[19]
port 11 nsew signal input
rlabel metal3 s 249200 19320 250000 19440 6 io_in[1]
port 12 nsew signal input
rlabel metal2 s 111522 249200 111578 250000 6 io_in[20]
port 13 nsew signal input
rlabel metal2 s 84750 249200 84806 250000 6 io_in[21]
port 14 nsew signal input
rlabel metal2 s 57978 249200 58034 250000 6 io_in[22]
port 15 nsew signal input
rlabel metal2 s 31206 249200 31262 250000 6 io_in[23]
port 16 nsew signal input
rlabel metal3 s 0 246984 800 247104 6 io_in[24]
port 17 nsew signal input
rlabel metal3 s 0 229848 800 229968 6 io_in[25]
port 18 nsew signal input
rlabel metal3 s 0 212848 800 212968 6 io_in[26]
port 19 nsew signal input
rlabel metal3 s 0 195848 800 195968 6 io_in[27]
port 20 nsew signal input
rlabel metal3 s 0 178712 800 178832 6 io_in[28]
port 21 nsew signal input
rlabel metal3 s 0 161712 800 161832 6 io_in[29]
port 22 nsew signal input
rlabel metal3 s 249200 36048 250000 36168 6 io_in[2]
port 23 nsew signal input
rlabel metal3 s 0 144712 800 144832 6 io_in[30]
port 24 nsew signal input
rlabel metal3 s 0 127712 800 127832 6 io_in[31]
port 25 nsew signal input
rlabel metal3 s 0 110576 800 110696 6 io_in[32]
port 26 nsew signal input
rlabel metal3 s 0 93576 800 93696 6 io_in[33]
port 27 nsew signal input
rlabel metal3 s 0 76576 800 76696 6 io_in[34]
port 28 nsew signal input
rlabel metal3 s 0 59440 800 59560 6 io_in[35]
port 29 nsew signal input
rlabel metal3 s 0 42440 800 42560 6 io_in[36]
port 30 nsew signal input
rlabel metal3 s 0 25440 800 25560 6 io_in[37]
port 31 nsew signal input
rlabel metal3 s 249200 52640 250000 52760 6 io_in[3]
port 32 nsew signal input
rlabel metal3 s 249200 69368 250000 69488 6 io_in[4]
port 33 nsew signal input
rlabel metal3 s 249200 85960 250000 86080 6 io_in[5]
port 34 nsew signal input
rlabel metal3 s 249200 102688 250000 102808 6 io_in[6]
port 35 nsew signal input
rlabel metal3 s 249200 119280 250000 119400 6 io_in[7]
port 36 nsew signal input
rlabel metal3 s 249200 136008 250000 136128 6 io_in[8]
port 37 nsew signal input
rlabel metal3 s 249200 152600 250000 152720 6 io_in[9]
port 38 nsew signal input
rlabel metal3 s 249200 13744 250000 13864 6 io_oeb[0]
port 39 nsew signal output
rlabel metal3 s 249200 180480 250000 180600 6 io_oeb[10]
port 40 nsew signal output
rlabel metal3 s 249200 197072 250000 197192 6 io_oeb[11]
port 41 nsew signal output
rlabel metal3 s 249200 213800 250000 213920 6 io_oeb[12]
port 42 nsew signal output
rlabel metal3 s 249200 230392 250000 230512 6 io_oeb[13]
port 43 nsew signal output
rlabel metal3 s 249200 247120 250000 247240 6 io_oeb[14]
port 44 nsew signal output
rlabel metal2 s 227534 249200 227590 250000 6 io_oeb[15]
port 45 nsew signal output
rlabel metal2 s 200762 249200 200818 250000 6 io_oeb[16]
port 46 nsew signal output
rlabel metal2 s 173990 249200 174046 250000 6 io_oeb[17]
port 47 nsew signal output
rlabel metal2 s 147218 249200 147274 250000 6 io_oeb[18]
port 48 nsew signal output
rlabel metal2 s 120446 249200 120502 250000 6 io_oeb[19]
port 49 nsew signal output
rlabel metal3 s 249200 30472 250000 30592 6 io_oeb[1]
port 50 nsew signal output
rlabel metal2 s 93674 249200 93730 250000 6 io_oeb[20]
port 51 nsew signal output
rlabel metal2 s 66902 249200 66958 250000 6 io_oeb[21]
port 52 nsew signal output
rlabel metal2 s 40130 249200 40186 250000 6 io_oeb[22]
port 53 nsew signal output
rlabel metal2 s 13358 249200 13414 250000 6 io_oeb[23]
port 54 nsew signal output
rlabel metal3 s 0 235560 800 235680 6 io_oeb[24]
port 55 nsew signal output
rlabel metal3 s 0 218560 800 218680 6 io_oeb[25]
port 56 nsew signal output
rlabel metal3 s 0 201560 800 201680 6 io_oeb[26]
port 57 nsew signal output
rlabel metal3 s 0 184424 800 184544 6 io_oeb[27]
port 58 nsew signal output
rlabel metal3 s 0 167424 800 167544 6 io_oeb[28]
port 59 nsew signal output
rlabel metal3 s 0 150424 800 150544 6 io_oeb[29]
port 60 nsew signal output
rlabel metal3 s 249200 47064 250000 47184 6 io_oeb[2]
port 61 nsew signal output
rlabel metal3 s 0 133288 800 133408 6 io_oeb[30]
port 62 nsew signal output
rlabel metal3 s 0 116288 800 116408 6 io_oeb[31]
port 63 nsew signal output
rlabel metal3 s 0 99288 800 99408 6 io_oeb[32]
port 64 nsew signal output
rlabel metal3 s 0 82152 800 82272 6 io_oeb[33]
port 65 nsew signal output
rlabel metal3 s 0 65152 800 65272 6 io_oeb[34]
port 66 nsew signal output
rlabel metal3 s 0 48152 800 48272 6 io_oeb[35]
port 67 nsew signal output
rlabel metal3 s 0 31016 800 31136 6 io_oeb[36]
port 68 nsew signal output
rlabel metal3 s 0 14016 800 14136 6 io_oeb[37]
port 69 nsew signal output
rlabel metal3 s 249200 63792 250000 63912 6 io_oeb[3]
port 70 nsew signal output
rlabel metal3 s 249200 80384 250000 80504 6 io_oeb[4]
port 71 nsew signal output
rlabel metal3 s 249200 97112 250000 97232 6 io_oeb[5]
port 72 nsew signal output
rlabel metal3 s 249200 113704 250000 113824 6 io_oeb[6]
port 73 nsew signal output
rlabel metal3 s 249200 130432 250000 130552 6 io_oeb[7]
port 74 nsew signal output
rlabel metal3 s 249200 147024 250000 147144 6 io_oeb[8]
port 75 nsew signal output
rlabel metal3 s 249200 163752 250000 163872 6 io_oeb[9]
port 76 nsew signal output
rlabel metal3 s 249200 8168 250000 8288 6 io_out[0]
port 77 nsew signal output
rlabel metal3 s 249200 174904 250000 175024 6 io_out[10]
port 78 nsew signal output
rlabel metal3 s 249200 191496 250000 191616 6 io_out[11]
port 79 nsew signal output
rlabel metal3 s 249200 208224 250000 208344 6 io_out[12]
port 80 nsew signal output
rlabel metal3 s 249200 224816 250000 224936 6 io_out[13]
port 81 nsew signal output
rlabel metal3 s 249200 241544 250000 241664 6 io_out[14]
port 82 nsew signal output
rlabel metal2 s 236458 249200 236514 250000 6 io_out[15]
port 83 nsew signal output
rlabel metal2 s 209686 249200 209742 250000 6 io_out[16]
port 84 nsew signal output
rlabel metal2 s 182914 249200 182970 250000 6 io_out[17]
port 85 nsew signal output
rlabel metal2 s 156142 249200 156198 250000 6 io_out[18]
port 86 nsew signal output
rlabel metal2 s 129370 249200 129426 250000 6 io_out[19]
port 87 nsew signal output
rlabel metal3 s 249200 24896 250000 25016 6 io_out[1]
port 88 nsew signal output
rlabel metal2 s 102598 249200 102654 250000 6 io_out[20]
port 89 nsew signal output
rlabel metal2 s 75826 249200 75882 250000 6 io_out[21]
port 90 nsew signal output
rlabel metal2 s 49054 249200 49110 250000 6 io_out[22]
port 91 nsew signal output
rlabel metal2 s 22282 249200 22338 250000 6 io_out[23]
port 92 nsew signal output
rlabel metal3 s 0 241272 800 241392 6 io_out[24]
port 93 nsew signal output
rlabel metal3 s 0 224272 800 224392 6 io_out[25]
port 94 nsew signal output
rlabel metal3 s 0 207136 800 207256 6 io_out[26]
port 95 nsew signal output
rlabel metal3 s 0 190136 800 190256 6 io_out[27]
port 96 nsew signal output
rlabel metal3 s 0 173136 800 173256 6 io_out[28]
port 97 nsew signal output
rlabel metal3 s 0 156000 800 156120 6 io_out[29]
port 98 nsew signal output
rlabel metal3 s 249200 41488 250000 41608 6 io_out[2]
port 99 nsew signal output
rlabel metal3 s 0 139000 800 139120 6 io_out[30]
port 100 nsew signal output
rlabel metal3 s 0 122000 800 122120 6 io_out[31]
port 101 nsew signal output
rlabel metal3 s 0 104864 800 104984 6 io_out[32]
port 102 nsew signal output
rlabel metal3 s 0 87864 800 87984 6 io_out[33]
port 103 nsew signal output
rlabel metal3 s 0 70864 800 70984 6 io_out[34]
port 104 nsew signal output
rlabel metal3 s 0 53728 800 53848 6 io_out[35]
port 105 nsew signal output
rlabel metal3 s 0 36728 800 36848 6 io_out[36]
port 106 nsew signal output
rlabel metal3 s 0 19728 800 19848 6 io_out[37]
port 107 nsew signal output
rlabel metal3 s 249200 58216 250000 58336 6 io_out[3]
port 108 nsew signal output
rlabel metal3 s 249200 74808 250000 74928 6 io_out[4]
port 109 nsew signal output
rlabel metal3 s 249200 91536 250000 91656 6 io_out[5]
port 110 nsew signal output
rlabel metal3 s 249200 108264 250000 108384 6 io_out[6]
port 111 nsew signal output
rlabel metal3 s 249200 124856 250000 124976 6 io_out[7]
port 112 nsew signal output
rlabel metal3 s 249200 141584 250000 141704 6 io_out[8]
port 113 nsew signal output
rlabel metal3 s 249200 158176 250000 158296 6 io_out[9]
port 114 nsew signal output
rlabel metal3 s 0 8304 800 8424 6 irq[0]
port 115 nsew signal output
rlabel metal2 s 4434 249200 4490 250000 6 irq[1]
port 116 nsew signal output
rlabel metal3 s 0 2728 800 2848 6 irq[2]
port 117 nsew signal output
rlabel metal2 s 54206 0 54262 800 6 la_data_in[0]
port 118 nsew signal input
rlabel metal2 s 207294 0 207350 800 6 la_data_in[100]
port 119 nsew signal input
rlabel metal2 s 208766 0 208822 800 6 la_data_in[101]
port 120 nsew signal input
rlabel metal2 s 210330 0 210386 800 6 la_data_in[102]
port 121 nsew signal input
rlabel metal2 s 211894 0 211950 800 6 la_data_in[103]
port 122 nsew signal input
rlabel metal2 s 213366 0 213422 800 6 la_data_in[104]
port 123 nsew signal input
rlabel metal2 s 214930 0 214986 800 6 la_data_in[105]
port 124 nsew signal input
rlabel metal2 s 216494 0 216550 800 6 la_data_in[106]
port 125 nsew signal input
rlabel metal2 s 217966 0 218022 800 6 la_data_in[107]
port 126 nsew signal input
rlabel metal2 s 219530 0 219586 800 6 la_data_in[108]
port 127 nsew signal input
rlabel metal2 s 221002 0 221058 800 6 la_data_in[109]
port 128 nsew signal input
rlabel metal2 s 69570 0 69626 800 6 la_data_in[10]
port 129 nsew signal input
rlabel metal2 s 222566 0 222622 800 6 la_data_in[110]
port 130 nsew signal input
rlabel metal2 s 224130 0 224186 800 6 la_data_in[111]
port 131 nsew signal input
rlabel metal2 s 225602 0 225658 800 6 la_data_in[112]
port 132 nsew signal input
rlabel metal2 s 227166 0 227222 800 6 la_data_in[113]
port 133 nsew signal input
rlabel metal2 s 228730 0 228786 800 6 la_data_in[114]
port 134 nsew signal input
rlabel metal2 s 230202 0 230258 800 6 la_data_in[115]
port 135 nsew signal input
rlabel metal2 s 231766 0 231822 800 6 la_data_in[116]
port 136 nsew signal input
rlabel metal2 s 233330 0 233386 800 6 la_data_in[117]
port 137 nsew signal input
rlabel metal2 s 234802 0 234858 800 6 la_data_in[118]
port 138 nsew signal input
rlabel metal2 s 236366 0 236422 800 6 la_data_in[119]
port 139 nsew signal input
rlabel metal2 s 71042 0 71098 800 6 la_data_in[11]
port 140 nsew signal input
rlabel metal2 s 237838 0 237894 800 6 la_data_in[120]
port 141 nsew signal input
rlabel metal2 s 239402 0 239458 800 6 la_data_in[121]
port 142 nsew signal input
rlabel metal2 s 240966 0 241022 800 6 la_data_in[122]
port 143 nsew signal input
rlabel metal2 s 242438 0 242494 800 6 la_data_in[123]
port 144 nsew signal input
rlabel metal2 s 244002 0 244058 800 6 la_data_in[124]
port 145 nsew signal input
rlabel metal2 s 245566 0 245622 800 6 la_data_in[125]
port 146 nsew signal input
rlabel metal2 s 247038 0 247094 800 6 la_data_in[126]
port 147 nsew signal input
rlabel metal2 s 248602 0 248658 800 6 la_data_in[127]
port 148 nsew signal input
rlabel metal2 s 72606 0 72662 800 6 la_data_in[12]
port 149 nsew signal input
rlabel metal2 s 74170 0 74226 800 6 la_data_in[13]
port 150 nsew signal input
rlabel metal2 s 75642 0 75698 800 6 la_data_in[14]
port 151 nsew signal input
rlabel metal2 s 77206 0 77262 800 6 la_data_in[15]
port 152 nsew signal input
rlabel metal2 s 78678 0 78734 800 6 la_data_in[16]
port 153 nsew signal input
rlabel metal2 s 80242 0 80298 800 6 la_data_in[17]
port 154 nsew signal input
rlabel metal2 s 81806 0 81862 800 6 la_data_in[18]
port 155 nsew signal input
rlabel metal2 s 83278 0 83334 800 6 la_data_in[19]
port 156 nsew signal input
rlabel metal2 s 55770 0 55826 800 6 la_data_in[1]
port 157 nsew signal input
rlabel metal2 s 84842 0 84898 800 6 la_data_in[20]
port 158 nsew signal input
rlabel metal2 s 86406 0 86462 800 6 la_data_in[21]
port 159 nsew signal input
rlabel metal2 s 87878 0 87934 800 6 la_data_in[22]
port 160 nsew signal input
rlabel metal2 s 89442 0 89498 800 6 la_data_in[23]
port 161 nsew signal input
rlabel metal2 s 90914 0 90970 800 6 la_data_in[24]
port 162 nsew signal input
rlabel metal2 s 92478 0 92534 800 6 la_data_in[25]
port 163 nsew signal input
rlabel metal2 s 94042 0 94098 800 6 la_data_in[26]
port 164 nsew signal input
rlabel metal2 s 95514 0 95570 800 6 la_data_in[27]
port 165 nsew signal input
rlabel metal2 s 97078 0 97134 800 6 la_data_in[28]
port 166 nsew signal input
rlabel metal2 s 98642 0 98698 800 6 la_data_in[29]
port 167 nsew signal input
rlabel metal2 s 57334 0 57390 800 6 la_data_in[2]
port 168 nsew signal input
rlabel metal2 s 100114 0 100170 800 6 la_data_in[30]
port 169 nsew signal input
rlabel metal2 s 101678 0 101734 800 6 la_data_in[31]
port 170 nsew signal input
rlabel metal2 s 103242 0 103298 800 6 la_data_in[32]
port 171 nsew signal input
rlabel metal2 s 104714 0 104770 800 6 la_data_in[33]
port 172 nsew signal input
rlabel metal2 s 106278 0 106334 800 6 la_data_in[34]
port 173 nsew signal input
rlabel metal2 s 107750 0 107806 800 6 la_data_in[35]
port 174 nsew signal input
rlabel metal2 s 109314 0 109370 800 6 la_data_in[36]
port 175 nsew signal input
rlabel metal2 s 110878 0 110934 800 6 la_data_in[37]
port 176 nsew signal input
rlabel metal2 s 112350 0 112406 800 6 la_data_in[38]
port 177 nsew signal input
rlabel metal2 s 113914 0 113970 800 6 la_data_in[39]
port 178 nsew signal input
rlabel metal2 s 58806 0 58862 800 6 la_data_in[3]
port 179 nsew signal input
rlabel metal2 s 115478 0 115534 800 6 la_data_in[40]
port 180 nsew signal input
rlabel metal2 s 116950 0 117006 800 6 la_data_in[41]
port 181 nsew signal input
rlabel metal2 s 118514 0 118570 800 6 la_data_in[42]
port 182 nsew signal input
rlabel metal2 s 120078 0 120134 800 6 la_data_in[43]
port 183 nsew signal input
rlabel metal2 s 121550 0 121606 800 6 la_data_in[44]
port 184 nsew signal input
rlabel metal2 s 123114 0 123170 800 6 la_data_in[45]
port 185 nsew signal input
rlabel metal2 s 124586 0 124642 800 6 la_data_in[46]
port 186 nsew signal input
rlabel metal2 s 126150 0 126206 800 6 la_data_in[47]
port 187 nsew signal input
rlabel metal2 s 127714 0 127770 800 6 la_data_in[48]
port 188 nsew signal input
rlabel metal2 s 129186 0 129242 800 6 la_data_in[49]
port 189 nsew signal input
rlabel metal2 s 60370 0 60426 800 6 la_data_in[4]
port 190 nsew signal input
rlabel metal2 s 130750 0 130806 800 6 la_data_in[50]
port 191 nsew signal input
rlabel metal2 s 132314 0 132370 800 6 la_data_in[51]
port 192 nsew signal input
rlabel metal2 s 133786 0 133842 800 6 la_data_in[52]
port 193 nsew signal input
rlabel metal2 s 135350 0 135406 800 6 la_data_in[53]
port 194 nsew signal input
rlabel metal2 s 136914 0 136970 800 6 la_data_in[54]
port 195 nsew signal input
rlabel metal2 s 138386 0 138442 800 6 la_data_in[55]
port 196 nsew signal input
rlabel metal2 s 139950 0 140006 800 6 la_data_in[56]
port 197 nsew signal input
rlabel metal2 s 141422 0 141478 800 6 la_data_in[57]
port 198 nsew signal input
rlabel metal2 s 142986 0 143042 800 6 la_data_in[58]
port 199 nsew signal input
rlabel metal2 s 144550 0 144606 800 6 la_data_in[59]
port 200 nsew signal input
rlabel metal2 s 61842 0 61898 800 6 la_data_in[5]
port 201 nsew signal input
rlabel metal2 s 146022 0 146078 800 6 la_data_in[60]
port 202 nsew signal input
rlabel metal2 s 147586 0 147642 800 6 la_data_in[61]
port 203 nsew signal input
rlabel metal2 s 149150 0 149206 800 6 la_data_in[62]
port 204 nsew signal input
rlabel metal2 s 150622 0 150678 800 6 la_data_in[63]
port 205 nsew signal input
rlabel metal2 s 152186 0 152242 800 6 la_data_in[64]
port 206 nsew signal input
rlabel metal2 s 153750 0 153806 800 6 la_data_in[65]
port 207 nsew signal input
rlabel metal2 s 155222 0 155278 800 6 la_data_in[66]
port 208 nsew signal input
rlabel metal2 s 156786 0 156842 800 6 la_data_in[67]
port 209 nsew signal input
rlabel metal2 s 158258 0 158314 800 6 la_data_in[68]
port 210 nsew signal input
rlabel metal2 s 159822 0 159878 800 6 la_data_in[69]
port 211 nsew signal input
rlabel metal2 s 63406 0 63462 800 6 la_data_in[6]
port 212 nsew signal input
rlabel metal2 s 161386 0 161442 800 6 la_data_in[70]
port 213 nsew signal input
rlabel metal2 s 162858 0 162914 800 6 la_data_in[71]
port 214 nsew signal input
rlabel metal2 s 164422 0 164478 800 6 la_data_in[72]
port 215 nsew signal input
rlabel metal2 s 165986 0 166042 800 6 la_data_in[73]
port 216 nsew signal input
rlabel metal2 s 167458 0 167514 800 6 la_data_in[74]
port 217 nsew signal input
rlabel metal2 s 169022 0 169078 800 6 la_data_in[75]
port 218 nsew signal input
rlabel metal2 s 170494 0 170550 800 6 la_data_in[76]
port 219 nsew signal input
rlabel metal2 s 172058 0 172114 800 6 la_data_in[77]
port 220 nsew signal input
rlabel metal2 s 173622 0 173678 800 6 la_data_in[78]
port 221 nsew signal input
rlabel metal2 s 175094 0 175150 800 6 la_data_in[79]
port 222 nsew signal input
rlabel metal2 s 64970 0 65026 800 6 la_data_in[7]
port 223 nsew signal input
rlabel metal2 s 176658 0 176714 800 6 la_data_in[80]
port 224 nsew signal input
rlabel metal2 s 178222 0 178278 800 6 la_data_in[81]
port 225 nsew signal input
rlabel metal2 s 179694 0 179750 800 6 la_data_in[82]
port 226 nsew signal input
rlabel metal2 s 181258 0 181314 800 6 la_data_in[83]
port 227 nsew signal input
rlabel metal2 s 182822 0 182878 800 6 la_data_in[84]
port 228 nsew signal input
rlabel metal2 s 184294 0 184350 800 6 la_data_in[85]
port 229 nsew signal input
rlabel metal2 s 185858 0 185914 800 6 la_data_in[86]
port 230 nsew signal input
rlabel metal2 s 187330 0 187386 800 6 la_data_in[87]
port 231 nsew signal input
rlabel metal2 s 188894 0 188950 800 6 la_data_in[88]
port 232 nsew signal input
rlabel metal2 s 190458 0 190514 800 6 la_data_in[89]
port 233 nsew signal input
rlabel metal2 s 66442 0 66498 800 6 la_data_in[8]
port 234 nsew signal input
rlabel metal2 s 191930 0 191986 800 6 la_data_in[90]
port 235 nsew signal input
rlabel metal2 s 193494 0 193550 800 6 la_data_in[91]
port 236 nsew signal input
rlabel metal2 s 195058 0 195114 800 6 la_data_in[92]
port 237 nsew signal input
rlabel metal2 s 196530 0 196586 800 6 la_data_in[93]
port 238 nsew signal input
rlabel metal2 s 198094 0 198150 800 6 la_data_in[94]
port 239 nsew signal input
rlabel metal2 s 199658 0 199714 800 6 la_data_in[95]
port 240 nsew signal input
rlabel metal2 s 201130 0 201186 800 6 la_data_in[96]
port 241 nsew signal input
rlabel metal2 s 202694 0 202750 800 6 la_data_in[97]
port 242 nsew signal input
rlabel metal2 s 204166 0 204222 800 6 la_data_in[98]
port 243 nsew signal input
rlabel metal2 s 205730 0 205786 800 6 la_data_in[99]
port 244 nsew signal input
rlabel metal2 s 68006 0 68062 800 6 la_data_in[9]
port 245 nsew signal input
rlabel metal2 s 54758 0 54814 800 6 la_data_out[0]
port 246 nsew signal output
rlabel metal2 s 207754 0 207810 800 6 la_data_out[100]
port 247 nsew signal output
rlabel metal2 s 209318 0 209374 800 6 la_data_out[101]
port 248 nsew signal output
rlabel metal2 s 210882 0 210938 800 6 la_data_out[102]
port 249 nsew signal output
rlabel metal2 s 212354 0 212410 800 6 la_data_out[103]
port 250 nsew signal output
rlabel metal2 s 213918 0 213974 800 6 la_data_out[104]
port 251 nsew signal output
rlabel metal2 s 215390 0 215446 800 6 la_data_out[105]
port 252 nsew signal output
rlabel metal2 s 216954 0 217010 800 6 la_data_out[106]
port 253 nsew signal output
rlabel metal2 s 218518 0 218574 800 6 la_data_out[107]
port 254 nsew signal output
rlabel metal2 s 219990 0 220046 800 6 la_data_out[108]
port 255 nsew signal output
rlabel metal2 s 221554 0 221610 800 6 la_data_out[109]
port 256 nsew signal output
rlabel metal2 s 70030 0 70086 800 6 la_data_out[10]
port 257 nsew signal output
rlabel metal2 s 223118 0 223174 800 6 la_data_out[110]
port 258 nsew signal output
rlabel metal2 s 224590 0 224646 800 6 la_data_out[111]
port 259 nsew signal output
rlabel metal2 s 226154 0 226210 800 6 la_data_out[112]
port 260 nsew signal output
rlabel metal2 s 227718 0 227774 800 6 la_data_out[113]
port 261 nsew signal output
rlabel metal2 s 229190 0 229246 800 6 la_data_out[114]
port 262 nsew signal output
rlabel metal2 s 230754 0 230810 800 6 la_data_out[115]
port 263 nsew signal output
rlabel metal2 s 232226 0 232282 800 6 la_data_out[116]
port 264 nsew signal output
rlabel metal2 s 233790 0 233846 800 6 la_data_out[117]
port 265 nsew signal output
rlabel metal2 s 235354 0 235410 800 6 la_data_out[118]
port 266 nsew signal output
rlabel metal2 s 236826 0 236882 800 6 la_data_out[119]
port 267 nsew signal output
rlabel metal2 s 71594 0 71650 800 6 la_data_out[11]
port 268 nsew signal output
rlabel metal2 s 238390 0 238446 800 6 la_data_out[120]
port 269 nsew signal output
rlabel metal2 s 239954 0 240010 800 6 la_data_out[121]
port 270 nsew signal output
rlabel metal2 s 241426 0 241482 800 6 la_data_out[122]
port 271 nsew signal output
rlabel metal2 s 242990 0 243046 800 6 la_data_out[123]
port 272 nsew signal output
rlabel metal2 s 244554 0 244610 800 6 la_data_out[124]
port 273 nsew signal output
rlabel metal2 s 246026 0 246082 800 6 la_data_out[125]
port 274 nsew signal output
rlabel metal2 s 247590 0 247646 800 6 la_data_out[126]
port 275 nsew signal output
rlabel metal2 s 249062 0 249118 800 6 la_data_out[127]
port 276 nsew signal output
rlabel metal2 s 73066 0 73122 800 6 la_data_out[12]
port 277 nsew signal output
rlabel metal2 s 74630 0 74686 800 6 la_data_out[13]
port 278 nsew signal output
rlabel metal2 s 76194 0 76250 800 6 la_data_out[14]
port 279 nsew signal output
rlabel metal2 s 77666 0 77722 800 6 la_data_out[15]
port 280 nsew signal output
rlabel metal2 s 79230 0 79286 800 6 la_data_out[16]
port 281 nsew signal output
rlabel metal2 s 80794 0 80850 800 6 la_data_out[17]
port 282 nsew signal output
rlabel metal2 s 82266 0 82322 800 6 la_data_out[18]
port 283 nsew signal output
rlabel metal2 s 83830 0 83886 800 6 la_data_out[19]
port 284 nsew signal output
rlabel metal2 s 56230 0 56286 800 6 la_data_out[1]
port 285 nsew signal output
rlabel metal2 s 85302 0 85358 800 6 la_data_out[20]
port 286 nsew signal output
rlabel metal2 s 86866 0 86922 800 6 la_data_out[21]
port 287 nsew signal output
rlabel metal2 s 88430 0 88486 800 6 la_data_out[22]
port 288 nsew signal output
rlabel metal2 s 89902 0 89958 800 6 la_data_out[23]
port 289 nsew signal output
rlabel metal2 s 91466 0 91522 800 6 la_data_out[24]
port 290 nsew signal output
rlabel metal2 s 93030 0 93086 800 6 la_data_out[25]
port 291 nsew signal output
rlabel metal2 s 94502 0 94558 800 6 la_data_out[26]
port 292 nsew signal output
rlabel metal2 s 96066 0 96122 800 6 la_data_out[27]
port 293 nsew signal output
rlabel metal2 s 97630 0 97686 800 6 la_data_out[28]
port 294 nsew signal output
rlabel metal2 s 99102 0 99158 800 6 la_data_out[29]
port 295 nsew signal output
rlabel metal2 s 57794 0 57850 800 6 la_data_out[2]
port 296 nsew signal output
rlabel metal2 s 100666 0 100722 800 6 la_data_out[30]
port 297 nsew signal output
rlabel metal2 s 102138 0 102194 800 6 la_data_out[31]
port 298 nsew signal output
rlabel metal2 s 103702 0 103758 800 6 la_data_out[32]
port 299 nsew signal output
rlabel metal2 s 105266 0 105322 800 6 la_data_out[33]
port 300 nsew signal output
rlabel metal2 s 106738 0 106794 800 6 la_data_out[34]
port 301 nsew signal output
rlabel metal2 s 108302 0 108358 800 6 la_data_out[35]
port 302 nsew signal output
rlabel metal2 s 109866 0 109922 800 6 la_data_out[36]
port 303 nsew signal output
rlabel metal2 s 111338 0 111394 800 6 la_data_out[37]
port 304 nsew signal output
rlabel metal2 s 112902 0 112958 800 6 la_data_out[38]
port 305 nsew signal output
rlabel metal2 s 114466 0 114522 800 6 la_data_out[39]
port 306 nsew signal output
rlabel metal2 s 59358 0 59414 800 6 la_data_out[3]
port 307 nsew signal output
rlabel metal2 s 115938 0 115994 800 6 la_data_out[40]
port 308 nsew signal output
rlabel metal2 s 117502 0 117558 800 6 la_data_out[41]
port 309 nsew signal output
rlabel metal2 s 118974 0 119030 800 6 la_data_out[42]
port 310 nsew signal output
rlabel metal2 s 120538 0 120594 800 6 la_data_out[43]
port 311 nsew signal output
rlabel metal2 s 122102 0 122158 800 6 la_data_out[44]
port 312 nsew signal output
rlabel metal2 s 123574 0 123630 800 6 la_data_out[45]
port 313 nsew signal output
rlabel metal2 s 125138 0 125194 800 6 la_data_out[46]
port 314 nsew signal output
rlabel metal2 s 126702 0 126758 800 6 la_data_out[47]
port 315 nsew signal output
rlabel metal2 s 128174 0 128230 800 6 la_data_out[48]
port 316 nsew signal output
rlabel metal2 s 129738 0 129794 800 6 la_data_out[49]
port 317 nsew signal output
rlabel metal2 s 60830 0 60886 800 6 la_data_out[4]
port 318 nsew signal output
rlabel metal2 s 131302 0 131358 800 6 la_data_out[50]
port 319 nsew signal output
rlabel metal2 s 132774 0 132830 800 6 la_data_out[51]
port 320 nsew signal output
rlabel metal2 s 134338 0 134394 800 6 la_data_out[52]
port 321 nsew signal output
rlabel metal2 s 135810 0 135866 800 6 la_data_out[53]
port 322 nsew signal output
rlabel metal2 s 137374 0 137430 800 6 la_data_out[54]
port 323 nsew signal output
rlabel metal2 s 138938 0 138994 800 6 la_data_out[55]
port 324 nsew signal output
rlabel metal2 s 140410 0 140466 800 6 la_data_out[56]
port 325 nsew signal output
rlabel metal2 s 141974 0 142030 800 6 la_data_out[57]
port 326 nsew signal output
rlabel metal2 s 143538 0 143594 800 6 la_data_out[58]
port 327 nsew signal output
rlabel metal2 s 145010 0 145066 800 6 la_data_out[59]
port 328 nsew signal output
rlabel metal2 s 62394 0 62450 800 6 la_data_out[5]
port 329 nsew signal output
rlabel metal2 s 146574 0 146630 800 6 la_data_out[60]
port 330 nsew signal output
rlabel metal2 s 148138 0 148194 800 6 la_data_out[61]
port 331 nsew signal output
rlabel metal2 s 149610 0 149666 800 6 la_data_out[62]
port 332 nsew signal output
rlabel metal2 s 151174 0 151230 800 6 la_data_out[63]
port 333 nsew signal output
rlabel metal2 s 152646 0 152702 800 6 la_data_out[64]
port 334 nsew signal output
rlabel metal2 s 154210 0 154266 800 6 la_data_out[65]
port 335 nsew signal output
rlabel metal2 s 155774 0 155830 800 6 la_data_out[66]
port 336 nsew signal output
rlabel metal2 s 157246 0 157302 800 6 la_data_out[67]
port 337 nsew signal output
rlabel metal2 s 158810 0 158866 800 6 la_data_out[68]
port 338 nsew signal output
rlabel metal2 s 160374 0 160430 800 6 la_data_out[69]
port 339 nsew signal output
rlabel metal2 s 63958 0 64014 800 6 la_data_out[6]
port 340 nsew signal output
rlabel metal2 s 161846 0 161902 800 6 la_data_out[70]
port 341 nsew signal output
rlabel metal2 s 163410 0 163466 800 6 la_data_out[71]
port 342 nsew signal output
rlabel metal2 s 164974 0 165030 800 6 la_data_out[72]
port 343 nsew signal output
rlabel metal2 s 166446 0 166502 800 6 la_data_out[73]
port 344 nsew signal output
rlabel metal2 s 168010 0 168066 800 6 la_data_out[74]
port 345 nsew signal output
rlabel metal2 s 169482 0 169538 800 6 la_data_out[75]
port 346 nsew signal output
rlabel metal2 s 171046 0 171102 800 6 la_data_out[76]
port 347 nsew signal output
rlabel metal2 s 172610 0 172666 800 6 la_data_out[77]
port 348 nsew signal output
rlabel metal2 s 174082 0 174138 800 6 la_data_out[78]
port 349 nsew signal output
rlabel metal2 s 175646 0 175702 800 6 la_data_out[79]
port 350 nsew signal output
rlabel metal2 s 65430 0 65486 800 6 la_data_out[7]
port 351 nsew signal output
rlabel metal2 s 177210 0 177266 800 6 la_data_out[80]
port 352 nsew signal output
rlabel metal2 s 178682 0 178738 800 6 la_data_out[81]
port 353 nsew signal output
rlabel metal2 s 180246 0 180302 800 6 la_data_out[82]
port 354 nsew signal output
rlabel metal2 s 181718 0 181774 800 6 la_data_out[83]
port 355 nsew signal output
rlabel metal2 s 183282 0 183338 800 6 la_data_out[84]
port 356 nsew signal output
rlabel metal2 s 184846 0 184902 800 6 la_data_out[85]
port 357 nsew signal output
rlabel metal2 s 186318 0 186374 800 6 la_data_out[86]
port 358 nsew signal output
rlabel metal2 s 187882 0 187938 800 6 la_data_out[87]
port 359 nsew signal output
rlabel metal2 s 189446 0 189502 800 6 la_data_out[88]
port 360 nsew signal output
rlabel metal2 s 190918 0 190974 800 6 la_data_out[89]
port 361 nsew signal output
rlabel metal2 s 66994 0 67050 800 6 la_data_out[8]
port 362 nsew signal output
rlabel metal2 s 192482 0 192538 800 6 la_data_out[90]
port 363 nsew signal output
rlabel metal2 s 194046 0 194102 800 6 la_data_out[91]
port 364 nsew signal output
rlabel metal2 s 195518 0 195574 800 6 la_data_out[92]
port 365 nsew signal output
rlabel metal2 s 197082 0 197138 800 6 la_data_out[93]
port 366 nsew signal output
rlabel metal2 s 198554 0 198610 800 6 la_data_out[94]
port 367 nsew signal output
rlabel metal2 s 200118 0 200174 800 6 la_data_out[95]
port 368 nsew signal output
rlabel metal2 s 201682 0 201738 800 6 la_data_out[96]
port 369 nsew signal output
rlabel metal2 s 203154 0 203210 800 6 la_data_out[97]
port 370 nsew signal output
rlabel metal2 s 204718 0 204774 800 6 la_data_out[98]
port 371 nsew signal output
rlabel metal2 s 206282 0 206338 800 6 la_data_out[99]
port 372 nsew signal output
rlabel metal2 s 68558 0 68614 800 6 la_data_out[9]
port 373 nsew signal output
rlabel metal2 s 55218 0 55274 800 6 la_oenb[0]
port 374 nsew signal input
rlabel metal2 s 208306 0 208362 800 6 la_oenb[100]
port 375 nsew signal input
rlabel metal2 s 209778 0 209834 800 6 la_oenb[101]
port 376 nsew signal input
rlabel metal2 s 211342 0 211398 800 6 la_oenb[102]
port 377 nsew signal input
rlabel metal2 s 212906 0 212962 800 6 la_oenb[103]
port 378 nsew signal input
rlabel metal2 s 214378 0 214434 800 6 la_oenb[104]
port 379 nsew signal input
rlabel metal2 s 215942 0 215998 800 6 la_oenb[105]
port 380 nsew signal input
rlabel metal2 s 217506 0 217562 800 6 la_oenb[106]
port 381 nsew signal input
rlabel metal2 s 218978 0 219034 800 6 la_oenb[107]
port 382 nsew signal input
rlabel metal2 s 220542 0 220598 800 6 la_oenb[108]
port 383 nsew signal input
rlabel metal2 s 222106 0 222162 800 6 la_oenb[109]
port 384 nsew signal input
rlabel metal2 s 70582 0 70638 800 6 la_oenb[10]
port 385 nsew signal input
rlabel metal2 s 223578 0 223634 800 6 la_oenb[110]
port 386 nsew signal input
rlabel metal2 s 225142 0 225198 800 6 la_oenb[111]
port 387 nsew signal input
rlabel metal2 s 226614 0 226670 800 6 la_oenb[112]
port 388 nsew signal input
rlabel metal2 s 228178 0 228234 800 6 la_oenb[113]
port 389 nsew signal input
rlabel metal2 s 229742 0 229798 800 6 la_oenb[114]
port 390 nsew signal input
rlabel metal2 s 231214 0 231270 800 6 la_oenb[115]
port 391 nsew signal input
rlabel metal2 s 232778 0 232834 800 6 la_oenb[116]
port 392 nsew signal input
rlabel metal2 s 234342 0 234398 800 6 la_oenb[117]
port 393 nsew signal input
rlabel metal2 s 235814 0 235870 800 6 la_oenb[118]
port 394 nsew signal input
rlabel metal2 s 237378 0 237434 800 6 la_oenb[119]
port 395 nsew signal input
rlabel metal2 s 72054 0 72110 800 6 la_oenb[11]
port 396 nsew signal input
rlabel metal2 s 238942 0 238998 800 6 la_oenb[120]
port 397 nsew signal input
rlabel metal2 s 240414 0 240470 800 6 la_oenb[121]
port 398 nsew signal input
rlabel metal2 s 241978 0 242034 800 6 la_oenb[122]
port 399 nsew signal input
rlabel metal2 s 243450 0 243506 800 6 la_oenb[123]
port 400 nsew signal input
rlabel metal2 s 245014 0 245070 800 6 la_oenb[124]
port 401 nsew signal input
rlabel metal2 s 246578 0 246634 800 6 la_oenb[125]
port 402 nsew signal input
rlabel metal2 s 248050 0 248106 800 6 la_oenb[126]
port 403 nsew signal input
rlabel metal2 s 249614 0 249670 800 6 la_oenb[127]
port 404 nsew signal input
rlabel metal2 s 73618 0 73674 800 6 la_oenb[12]
port 405 nsew signal input
rlabel metal2 s 75182 0 75238 800 6 la_oenb[13]
port 406 nsew signal input
rlabel metal2 s 76654 0 76710 800 6 la_oenb[14]
port 407 nsew signal input
rlabel metal2 s 78218 0 78274 800 6 la_oenb[15]
port 408 nsew signal input
rlabel metal2 s 79782 0 79838 800 6 la_oenb[16]
port 409 nsew signal input
rlabel metal2 s 81254 0 81310 800 6 la_oenb[17]
port 410 nsew signal input
rlabel metal2 s 82818 0 82874 800 6 la_oenb[18]
port 411 nsew signal input
rlabel metal2 s 84290 0 84346 800 6 la_oenb[19]
port 412 nsew signal input
rlabel metal2 s 56782 0 56838 800 6 la_oenb[1]
port 413 nsew signal input
rlabel metal2 s 85854 0 85910 800 6 la_oenb[20]
port 414 nsew signal input
rlabel metal2 s 87418 0 87474 800 6 la_oenb[21]
port 415 nsew signal input
rlabel metal2 s 88890 0 88946 800 6 la_oenb[22]
port 416 nsew signal input
rlabel metal2 s 90454 0 90510 800 6 la_oenb[23]
port 417 nsew signal input
rlabel metal2 s 92018 0 92074 800 6 la_oenb[24]
port 418 nsew signal input
rlabel metal2 s 93490 0 93546 800 6 la_oenb[25]
port 419 nsew signal input
rlabel metal2 s 95054 0 95110 800 6 la_oenb[26]
port 420 nsew signal input
rlabel metal2 s 96526 0 96582 800 6 la_oenb[27]
port 421 nsew signal input
rlabel metal2 s 98090 0 98146 800 6 la_oenb[28]
port 422 nsew signal input
rlabel metal2 s 99654 0 99710 800 6 la_oenb[29]
port 423 nsew signal input
rlabel metal2 s 58346 0 58402 800 6 la_oenb[2]
port 424 nsew signal input
rlabel metal2 s 101126 0 101182 800 6 la_oenb[30]
port 425 nsew signal input
rlabel metal2 s 102690 0 102746 800 6 la_oenb[31]
port 426 nsew signal input
rlabel metal2 s 104254 0 104310 800 6 la_oenb[32]
port 427 nsew signal input
rlabel metal2 s 105726 0 105782 800 6 la_oenb[33]
port 428 nsew signal input
rlabel metal2 s 107290 0 107346 800 6 la_oenb[34]
port 429 nsew signal input
rlabel metal2 s 108854 0 108910 800 6 la_oenb[35]
port 430 nsew signal input
rlabel metal2 s 110326 0 110382 800 6 la_oenb[36]
port 431 nsew signal input
rlabel metal2 s 111890 0 111946 800 6 la_oenb[37]
port 432 nsew signal input
rlabel metal2 s 113362 0 113418 800 6 la_oenb[38]
port 433 nsew signal input
rlabel metal2 s 114926 0 114982 800 6 la_oenb[39]
port 434 nsew signal input
rlabel metal2 s 59818 0 59874 800 6 la_oenb[3]
port 435 nsew signal input
rlabel metal2 s 116490 0 116546 800 6 la_oenb[40]
port 436 nsew signal input
rlabel metal2 s 117962 0 118018 800 6 la_oenb[41]
port 437 nsew signal input
rlabel metal2 s 119526 0 119582 800 6 la_oenb[42]
port 438 nsew signal input
rlabel metal2 s 121090 0 121146 800 6 la_oenb[43]
port 439 nsew signal input
rlabel metal2 s 122562 0 122618 800 6 la_oenb[44]
port 440 nsew signal input
rlabel metal2 s 124126 0 124182 800 6 la_oenb[45]
port 441 nsew signal input
rlabel metal2 s 125690 0 125746 800 6 la_oenb[46]
port 442 nsew signal input
rlabel metal2 s 127162 0 127218 800 6 la_oenb[47]
port 443 nsew signal input
rlabel metal2 s 128726 0 128782 800 6 la_oenb[48]
port 444 nsew signal input
rlabel metal2 s 130198 0 130254 800 6 la_oenb[49]
port 445 nsew signal input
rlabel metal2 s 61382 0 61438 800 6 la_oenb[4]
port 446 nsew signal input
rlabel metal2 s 131762 0 131818 800 6 la_oenb[50]
port 447 nsew signal input
rlabel metal2 s 133326 0 133382 800 6 la_oenb[51]
port 448 nsew signal input
rlabel metal2 s 134798 0 134854 800 6 la_oenb[52]
port 449 nsew signal input
rlabel metal2 s 136362 0 136418 800 6 la_oenb[53]
port 450 nsew signal input
rlabel metal2 s 137926 0 137982 800 6 la_oenb[54]
port 451 nsew signal input
rlabel metal2 s 139398 0 139454 800 6 la_oenb[55]
port 452 nsew signal input
rlabel metal2 s 140962 0 141018 800 6 la_oenb[56]
port 453 nsew signal input
rlabel metal2 s 142526 0 142582 800 6 la_oenb[57]
port 454 nsew signal input
rlabel metal2 s 143998 0 144054 800 6 la_oenb[58]
port 455 nsew signal input
rlabel metal2 s 145562 0 145618 800 6 la_oenb[59]
port 456 nsew signal input
rlabel metal2 s 62946 0 63002 800 6 la_oenb[5]
port 457 nsew signal input
rlabel metal2 s 147034 0 147090 800 6 la_oenb[60]
port 458 nsew signal input
rlabel metal2 s 148598 0 148654 800 6 la_oenb[61]
port 459 nsew signal input
rlabel metal2 s 150162 0 150218 800 6 la_oenb[62]
port 460 nsew signal input
rlabel metal2 s 151634 0 151690 800 6 la_oenb[63]
port 461 nsew signal input
rlabel metal2 s 153198 0 153254 800 6 la_oenb[64]
port 462 nsew signal input
rlabel metal2 s 154762 0 154818 800 6 la_oenb[65]
port 463 nsew signal input
rlabel metal2 s 156234 0 156290 800 6 la_oenb[66]
port 464 nsew signal input
rlabel metal2 s 157798 0 157854 800 6 la_oenb[67]
port 465 nsew signal input
rlabel metal2 s 159362 0 159418 800 6 la_oenb[68]
port 466 nsew signal input
rlabel metal2 s 160834 0 160890 800 6 la_oenb[69]
port 467 nsew signal input
rlabel metal2 s 64418 0 64474 800 6 la_oenb[6]
port 468 nsew signal input
rlabel metal2 s 162398 0 162454 800 6 la_oenb[70]
port 469 nsew signal input
rlabel metal2 s 163870 0 163926 800 6 la_oenb[71]
port 470 nsew signal input
rlabel metal2 s 165434 0 165490 800 6 la_oenb[72]
port 471 nsew signal input
rlabel metal2 s 166998 0 167054 800 6 la_oenb[73]
port 472 nsew signal input
rlabel metal2 s 168470 0 168526 800 6 la_oenb[74]
port 473 nsew signal input
rlabel metal2 s 170034 0 170090 800 6 la_oenb[75]
port 474 nsew signal input
rlabel metal2 s 171598 0 171654 800 6 la_oenb[76]
port 475 nsew signal input
rlabel metal2 s 173070 0 173126 800 6 la_oenb[77]
port 476 nsew signal input
rlabel metal2 s 174634 0 174690 800 6 la_oenb[78]
port 477 nsew signal input
rlabel metal2 s 176106 0 176162 800 6 la_oenb[79]
port 478 nsew signal input
rlabel metal2 s 65982 0 66038 800 6 la_oenb[7]
port 479 nsew signal input
rlabel metal2 s 177670 0 177726 800 6 la_oenb[80]
port 480 nsew signal input
rlabel metal2 s 179234 0 179290 800 6 la_oenb[81]
port 481 nsew signal input
rlabel metal2 s 180706 0 180762 800 6 la_oenb[82]
port 482 nsew signal input
rlabel metal2 s 182270 0 182326 800 6 la_oenb[83]
port 483 nsew signal input
rlabel metal2 s 183834 0 183890 800 6 la_oenb[84]
port 484 nsew signal input
rlabel metal2 s 185306 0 185362 800 6 la_oenb[85]
port 485 nsew signal input
rlabel metal2 s 186870 0 186926 800 6 la_oenb[86]
port 486 nsew signal input
rlabel metal2 s 188434 0 188490 800 6 la_oenb[87]
port 487 nsew signal input
rlabel metal2 s 189906 0 189962 800 6 la_oenb[88]
port 488 nsew signal input
rlabel metal2 s 191470 0 191526 800 6 la_oenb[89]
port 489 nsew signal input
rlabel metal2 s 67454 0 67510 800 6 la_oenb[8]
port 490 nsew signal input
rlabel metal2 s 192942 0 192998 800 6 la_oenb[90]
port 491 nsew signal input
rlabel metal2 s 194506 0 194562 800 6 la_oenb[91]
port 492 nsew signal input
rlabel metal2 s 196070 0 196126 800 6 la_oenb[92]
port 493 nsew signal input
rlabel metal2 s 197542 0 197598 800 6 la_oenb[93]
port 494 nsew signal input
rlabel metal2 s 199106 0 199162 800 6 la_oenb[94]
port 495 nsew signal input
rlabel metal2 s 200670 0 200726 800 6 la_oenb[95]
port 496 nsew signal input
rlabel metal2 s 202142 0 202198 800 6 la_oenb[96]
port 497 nsew signal input
rlabel metal2 s 203706 0 203762 800 6 la_oenb[97]
port 498 nsew signal input
rlabel metal2 s 205270 0 205326 800 6 la_oenb[98]
port 499 nsew signal input
rlabel metal2 s 206742 0 206798 800 6 la_oenb[99]
port 500 nsew signal input
rlabel metal2 s 69018 0 69074 800 6 la_oenb[9]
port 501 nsew signal input
rlabel metal4 s 4208 2128 4528 247568 6 vccd1
port 502 nsew power input
rlabel metal4 s 34928 2128 35248 247568 6 vccd1
port 502 nsew power input
rlabel metal4 s 65648 2128 65968 247568 6 vccd1
port 502 nsew power input
rlabel metal4 s 96368 2128 96688 247568 6 vccd1
port 502 nsew power input
rlabel metal4 s 127088 2128 127408 247568 6 vccd1
port 502 nsew power input
rlabel metal4 s 157808 2128 158128 247568 6 vccd1
port 502 nsew power input
rlabel metal4 s 188528 2128 188848 247568 6 vccd1
port 502 nsew power input
rlabel metal4 s 219248 2128 219568 247568 6 vccd1
port 502 nsew power input
rlabel metal4 s 19568 2128 19888 247568 6 vssd1
port 503 nsew ground input
rlabel metal4 s 50288 2128 50608 247568 6 vssd1
port 503 nsew ground input
rlabel metal4 s 81008 2128 81328 247568 6 vssd1
port 503 nsew ground input
rlabel metal4 s 111728 2128 112048 247568 6 vssd1
port 503 nsew ground input
rlabel metal4 s 142448 2128 142768 247568 6 vssd1
port 503 nsew ground input
rlabel metal4 s 173168 2128 173488 247568 6 vssd1
port 503 nsew ground input
rlabel metal4 s 203888 2128 204208 247568 6 vssd1
port 503 nsew ground input
rlabel metal4 s 234608 2128 234928 247568 6 vssd1
port 503 nsew ground input
rlabel metal2 s 202 0 258 800 6 wb_clk_i
port 504 nsew signal input
rlabel metal2 s 662 0 718 800 6 wb_rst_i
port 505 nsew signal input
rlabel metal2 s 1214 0 1270 800 6 wbs_ack_o
port 506 nsew signal output
rlabel metal2 s 3238 0 3294 800 6 wbs_adr_i[0]
port 507 nsew signal input
rlabel metal2 s 20534 0 20590 800 6 wbs_adr_i[10]
port 508 nsew signal input
rlabel metal2 s 22098 0 22154 800 6 wbs_adr_i[11]
port 509 nsew signal input
rlabel metal2 s 23662 0 23718 800 6 wbs_adr_i[12]
port 510 nsew signal input
rlabel metal2 s 25134 0 25190 800 6 wbs_adr_i[13]
port 511 nsew signal input
rlabel metal2 s 26698 0 26754 800 6 wbs_adr_i[14]
port 512 nsew signal input
rlabel metal2 s 28170 0 28226 800 6 wbs_adr_i[15]
port 513 nsew signal input
rlabel metal2 s 29734 0 29790 800 6 wbs_adr_i[16]
port 514 nsew signal input
rlabel metal2 s 31298 0 31354 800 6 wbs_adr_i[17]
port 515 nsew signal input
rlabel metal2 s 32770 0 32826 800 6 wbs_adr_i[18]
port 516 nsew signal input
rlabel metal2 s 34334 0 34390 800 6 wbs_adr_i[19]
port 517 nsew signal input
rlabel metal2 s 5262 0 5318 800 6 wbs_adr_i[1]
port 518 nsew signal input
rlabel metal2 s 35898 0 35954 800 6 wbs_adr_i[20]
port 519 nsew signal input
rlabel metal2 s 37370 0 37426 800 6 wbs_adr_i[21]
port 520 nsew signal input
rlabel metal2 s 38934 0 38990 800 6 wbs_adr_i[22]
port 521 nsew signal input
rlabel metal2 s 40498 0 40554 800 6 wbs_adr_i[23]
port 522 nsew signal input
rlabel metal2 s 41970 0 42026 800 6 wbs_adr_i[24]
port 523 nsew signal input
rlabel metal2 s 43534 0 43590 800 6 wbs_adr_i[25]
port 524 nsew signal input
rlabel metal2 s 45006 0 45062 800 6 wbs_adr_i[26]
port 525 nsew signal input
rlabel metal2 s 46570 0 46626 800 6 wbs_adr_i[27]
port 526 nsew signal input
rlabel metal2 s 48134 0 48190 800 6 wbs_adr_i[28]
port 527 nsew signal input
rlabel metal2 s 49606 0 49662 800 6 wbs_adr_i[29]
port 528 nsew signal input
rlabel metal2 s 7286 0 7342 800 6 wbs_adr_i[2]
port 529 nsew signal input
rlabel metal2 s 51170 0 51226 800 6 wbs_adr_i[30]
port 530 nsew signal input
rlabel metal2 s 52734 0 52790 800 6 wbs_adr_i[31]
port 531 nsew signal input
rlabel metal2 s 9310 0 9366 800 6 wbs_adr_i[3]
port 532 nsew signal input
rlabel metal2 s 11334 0 11390 800 6 wbs_adr_i[4]
port 533 nsew signal input
rlabel metal2 s 12898 0 12954 800 6 wbs_adr_i[5]
port 534 nsew signal input
rlabel metal2 s 14462 0 14518 800 6 wbs_adr_i[6]
port 535 nsew signal input
rlabel metal2 s 15934 0 15990 800 6 wbs_adr_i[7]
port 536 nsew signal input
rlabel metal2 s 17498 0 17554 800 6 wbs_adr_i[8]
port 537 nsew signal input
rlabel metal2 s 19062 0 19118 800 6 wbs_adr_i[9]
port 538 nsew signal input
rlabel metal2 s 1674 0 1730 800 6 wbs_cyc_i
port 539 nsew signal input
rlabel metal2 s 3698 0 3754 800 6 wbs_dat_i[0]
port 540 nsew signal input
rlabel metal2 s 21086 0 21142 800 6 wbs_dat_i[10]
port 541 nsew signal input
rlabel metal2 s 22558 0 22614 800 6 wbs_dat_i[11]
port 542 nsew signal input
rlabel metal2 s 24122 0 24178 800 6 wbs_dat_i[12]
port 543 nsew signal input
rlabel metal2 s 25686 0 25742 800 6 wbs_dat_i[13]
port 544 nsew signal input
rlabel metal2 s 27158 0 27214 800 6 wbs_dat_i[14]
port 545 nsew signal input
rlabel metal2 s 28722 0 28778 800 6 wbs_dat_i[15]
port 546 nsew signal input
rlabel metal2 s 30286 0 30342 800 6 wbs_dat_i[16]
port 547 nsew signal input
rlabel metal2 s 31758 0 31814 800 6 wbs_dat_i[17]
port 548 nsew signal input
rlabel metal2 s 33322 0 33378 800 6 wbs_dat_i[18]
port 549 nsew signal input
rlabel metal2 s 34886 0 34942 800 6 wbs_dat_i[19]
port 550 nsew signal input
rlabel metal2 s 5722 0 5778 800 6 wbs_dat_i[1]
port 551 nsew signal input
rlabel metal2 s 36358 0 36414 800 6 wbs_dat_i[20]
port 552 nsew signal input
rlabel metal2 s 37922 0 37978 800 6 wbs_dat_i[21]
port 553 nsew signal input
rlabel metal2 s 39394 0 39450 800 6 wbs_dat_i[22]
port 554 nsew signal input
rlabel metal2 s 40958 0 41014 800 6 wbs_dat_i[23]
port 555 nsew signal input
rlabel metal2 s 42522 0 42578 800 6 wbs_dat_i[24]
port 556 nsew signal input
rlabel metal2 s 43994 0 44050 800 6 wbs_dat_i[25]
port 557 nsew signal input
rlabel metal2 s 45558 0 45614 800 6 wbs_dat_i[26]
port 558 nsew signal input
rlabel metal2 s 47122 0 47178 800 6 wbs_dat_i[27]
port 559 nsew signal input
rlabel metal2 s 48594 0 48650 800 6 wbs_dat_i[28]
port 560 nsew signal input
rlabel metal2 s 50158 0 50214 800 6 wbs_dat_i[29]
port 561 nsew signal input
rlabel metal2 s 7838 0 7894 800 6 wbs_dat_i[2]
port 562 nsew signal input
rlabel metal2 s 51722 0 51778 800 6 wbs_dat_i[30]
port 563 nsew signal input
rlabel metal2 s 53194 0 53250 800 6 wbs_dat_i[31]
port 564 nsew signal input
rlabel metal2 s 9862 0 9918 800 6 wbs_dat_i[3]
port 565 nsew signal input
rlabel metal2 s 11886 0 11942 800 6 wbs_dat_i[4]
port 566 nsew signal input
rlabel metal2 s 13450 0 13506 800 6 wbs_dat_i[5]
port 567 nsew signal input
rlabel metal2 s 14922 0 14978 800 6 wbs_dat_i[6]
port 568 nsew signal input
rlabel metal2 s 16486 0 16542 800 6 wbs_dat_i[7]
port 569 nsew signal input
rlabel metal2 s 18050 0 18106 800 6 wbs_dat_i[8]
port 570 nsew signal input
rlabel metal2 s 19522 0 19578 800 6 wbs_dat_i[9]
port 571 nsew signal input
rlabel metal2 s 4250 0 4306 800 6 wbs_dat_o[0]
port 572 nsew signal output
rlabel metal2 s 21546 0 21602 800 6 wbs_dat_o[10]
port 573 nsew signal output
rlabel metal2 s 23110 0 23166 800 6 wbs_dat_o[11]
port 574 nsew signal output
rlabel metal2 s 24674 0 24730 800 6 wbs_dat_o[12]
port 575 nsew signal output
rlabel metal2 s 26146 0 26202 800 6 wbs_dat_o[13]
port 576 nsew signal output
rlabel metal2 s 27710 0 27766 800 6 wbs_dat_o[14]
port 577 nsew signal output
rlabel metal2 s 29274 0 29330 800 6 wbs_dat_o[15]
port 578 nsew signal output
rlabel metal2 s 30746 0 30802 800 6 wbs_dat_o[16]
port 579 nsew signal output
rlabel metal2 s 32310 0 32366 800 6 wbs_dat_o[17]
port 580 nsew signal output
rlabel metal2 s 33782 0 33838 800 6 wbs_dat_o[18]
port 581 nsew signal output
rlabel metal2 s 35346 0 35402 800 6 wbs_dat_o[19]
port 582 nsew signal output
rlabel metal2 s 6274 0 6330 800 6 wbs_dat_o[1]
port 583 nsew signal output
rlabel metal2 s 36910 0 36966 800 6 wbs_dat_o[20]
port 584 nsew signal output
rlabel metal2 s 38382 0 38438 800 6 wbs_dat_o[21]
port 585 nsew signal output
rlabel metal2 s 39946 0 40002 800 6 wbs_dat_o[22]
port 586 nsew signal output
rlabel metal2 s 41510 0 41566 800 6 wbs_dat_o[23]
port 587 nsew signal output
rlabel metal2 s 42982 0 43038 800 6 wbs_dat_o[24]
port 588 nsew signal output
rlabel metal2 s 44546 0 44602 800 6 wbs_dat_o[25]
port 589 nsew signal output
rlabel metal2 s 46110 0 46166 800 6 wbs_dat_o[26]
port 590 nsew signal output
rlabel metal2 s 47582 0 47638 800 6 wbs_dat_o[27]
port 591 nsew signal output
rlabel metal2 s 49146 0 49202 800 6 wbs_dat_o[28]
port 592 nsew signal output
rlabel metal2 s 50618 0 50674 800 6 wbs_dat_o[29]
port 593 nsew signal output
rlabel metal2 s 8298 0 8354 800 6 wbs_dat_o[2]
port 594 nsew signal output
rlabel metal2 s 52182 0 52238 800 6 wbs_dat_o[30]
port 595 nsew signal output
rlabel metal2 s 53746 0 53802 800 6 wbs_dat_o[31]
port 596 nsew signal output
rlabel metal2 s 10322 0 10378 800 6 wbs_dat_o[3]
port 597 nsew signal output
rlabel metal2 s 12438 0 12494 800 6 wbs_dat_o[4]
port 598 nsew signal output
rlabel metal2 s 13910 0 13966 800 6 wbs_dat_o[5]
port 599 nsew signal output
rlabel metal2 s 15474 0 15530 800 6 wbs_dat_o[6]
port 600 nsew signal output
rlabel metal2 s 16946 0 17002 800 6 wbs_dat_o[7]
port 601 nsew signal output
rlabel metal2 s 18510 0 18566 800 6 wbs_dat_o[8]
port 602 nsew signal output
rlabel metal2 s 20074 0 20130 800 6 wbs_dat_o[9]
port 603 nsew signal output
rlabel metal2 s 4710 0 4766 800 6 wbs_sel_i[0]
port 604 nsew signal input
rlabel metal2 s 6826 0 6882 800 6 wbs_sel_i[1]
port 605 nsew signal input
rlabel metal2 s 8850 0 8906 800 6 wbs_sel_i[2]
port 606 nsew signal input
rlabel metal2 s 10874 0 10930 800 6 wbs_sel_i[3]
port 607 nsew signal input
rlabel metal2 s 2226 0 2282 800 6 wbs_stb_i
port 608 nsew signal input
rlabel metal2 s 2686 0 2742 800 6 wbs_we_i
port 609 nsew signal input
<< properties >>
string FIXED_BBOX 0 0 250000 250000
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 44443362
string GDS_FILE /home/fatihgulakar/638_proje/shooting_game_verilog/openlane/user_proj_example/runs/user_proj_example/results/finishing/user_proj_example.magic.gds
string GDS_START 1775670
<< end >>

