module obj_p(
    input [5:0]  x,
    input [5:0]  y,
    input [3:0]  dir,
    input        en,
    output [1:0] data
);
    wire [1:0] rom [0:3][0:39][0:39] = { 
	 { { 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b10 , 2'b10 , 2'b10 , 2'b10 , 2'b10 , 2'b10 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 },
		{ 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b10 , 2'b10 , 2'b11 , 2'b11 , 2'b10 , 2'b10 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 },
		{ 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b10 , 2'b11 , 2'b11 , 2'b10 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 },
		{ 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b10 , 2'b11 , 2'b11 , 2'b10 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 },
		{ 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b10 , 2'b11 , 2'b11 , 2'b10 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 },
		{ 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b10 , 2'b11 , 2'b11 , 2'b10 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 },
		{ 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b10 , 2'b10 , 2'b10 , 2'b10 , 2'b10 , 2'b10 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b10 , 2'b11 , 2'b11 , 2'b10 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 },
		{ 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b10 , 2'b10 , 2'b10 , 2'b10 , 2'b10 , 2'b10 , 2'b00 , 2'b00 , 2'b00 , 2'b10 , 2'b10 , 2'b11 , 2'b11 , 2'b11 , 2'b11 , 2'b10 , 2'b10 , 2'b00 , 2'b00 , 2'b00 , 2'b10 , 2'b11 , 2'b11 , 2'b10 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 },
		{ 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b10 , 2'b10 , 2'b11 , 2'b11 , 2'b11 , 2'b11 , 2'b10 , 2'b10 , 2'b00 , 2'b00 , 2'b10 , 2'b11 , 2'b11 , 2'b11 , 2'b11 , 2'b11 , 2'b11 , 2'b10 , 2'b10 , 2'b00 , 2'b00 , 2'b10 , 2'b11 , 2'b11 , 2'b10 , 2'b10 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 },
		{ 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b10 , 2'b10 , 2'b11 , 2'b11 , 2'b11 , 2'b11 , 2'b11 , 2'b11 , 2'b10 , 2'b10 , 2'b00 , 2'b10 , 2'b11 , 2'b11 , 2'b11 , 2'b11 , 2'b11 , 2'b11 , 2'b11 , 2'b10 , 2'b00 , 2'b00 , 2'b10 , 2'b11 , 2'b11 , 2'b10 , 2'b10 , 2'b10 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 },
		{ 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b10 , 2'b11 , 2'b11 , 2'b11 , 2'b11 , 2'b11 , 2'b11 , 2'b10 , 2'b10 , 2'b10 , 2'b10 , 2'b10 , 2'b10 , 2'b10 , 2'b10 , 2'b10 , 2'b10 , 2'b10 , 2'b10 , 2'b10 , 2'b00 , 2'b00 , 2'b10 , 2'b11 , 2'b11 , 2'b10 , 2'b01 , 2'b10 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 },
		{ 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b10 , 2'b11 , 2'b11 , 2'b11 , 2'b11 , 2'b10 , 2'b10 , 2'b10 , 2'b10 , 2'b10 , 2'b10 , 2'b10 , 2'b10 , 2'b10 , 2'b10 , 2'b10 , 2'b10 , 2'b10 , 2'b10 , 2'b10 , 2'b10 , 2'b00 , 2'b10 , 2'b11 , 2'b11 , 2'b10 , 2'b01 , 2'b10 , 2'b10 , 2'b10 , 2'b10 , 2'b10 , 2'b10 },
		{ 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b10 , 2'b11 , 2'b11 , 2'b11 , 2'b11 , 2'b10 , 2'b10 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b10 , 2'b10 , 2'b00 , 2'b10 , 2'b11 , 2'b11 , 2'b10 , 2'b01 , 2'b01 , 2'b10 , 2'b10 , 2'b11 , 2'b11 , 2'b10 },
		{ 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b10 , 2'b11 , 2'b11 , 2'b10 , 2'b10 , 2'b10 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b10 , 2'b10 , 2'b10 , 2'b11 , 2'b11 , 2'b10 , 2'b01 , 2'b01 , 2'b01 , 2'b10 , 2'b11 , 2'b11 , 2'b10 },
		{ 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b10 , 2'b11 , 2'b10 , 2'b10 , 2'b10 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b10 , 2'b10 , 2'b11 , 2'b11 , 2'b10 , 2'b10 , 2'b01 , 2'b01 , 2'b10 , 2'b10 , 2'b11 , 2'b10 },
		{ 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b10 , 2'b10 , 2'b10 , 2'b10 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b10 , 2'b10 , 2'b11 , 2'b10 , 2'b10 , 2'b01 , 2'b01 , 2'b01 , 2'b10 , 2'b10 , 2'b10 },
		{ 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b10 , 2'b10 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b10 , 2'b10 , 2'b10 , 2'b10 , 2'b01 , 2'b01 , 2'b01 , 2'b10 , 2'b00 , 2'b00 },
		{ 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b10 , 2'b10 , 2'b10 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b10 , 2'b10 , 2'b10 , 2'b01 , 2'b01 , 2'b01 , 2'b10 , 2'b00 , 2'b00 },
		{ 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b10 , 2'b10 , 2'b10 , 2'b10 , 2'b10 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b10 , 2'b10 , 2'b10 , 2'b01 , 2'b01 , 2'b01 , 2'b10 , 2'b00 , 2'b00 },
		{ 2'b00 , 2'b00 , 2'b10 , 2'b10 , 2'b10 , 2'b01 , 2'b10 , 2'b10 , 2'b10 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b10 , 2'b10 , 2'b10 , 2'b01 , 2'b01 , 2'b01 , 2'b10 , 2'b00 , 2'b00 },
		{ 2'b00 , 2'b00 , 2'b10 , 2'b10 , 2'b01 , 2'b01 , 2'b10 , 2'b10 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b10 , 2'b10 , 2'b01 , 2'b01 , 2'b01 , 2'b10 , 2'b00 , 2'b00 },
		{ 2'b00 , 2'b00 , 2'b10 , 2'b01 , 2'b01 , 2'b01 , 2'b10 , 2'b10 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b10 , 2'b10 , 2'b01 , 2'b01 , 2'b01 , 2'b10 , 2'b00 , 2'b00 },
		{ 2'b00 , 2'b00 , 2'b10 , 2'b01 , 2'b01 , 2'b01 , 2'b10 , 2'b10 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b10 , 2'b10 , 2'b10 , 2'b01 , 2'b01 , 2'b01 , 2'b10 , 2'b00 , 2'b00 },
		{ 2'b00 , 2'b00 , 2'b10 , 2'b01 , 2'b01 , 2'b01 , 2'b10 , 2'b10 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b10 , 2'b10 , 2'b01 , 2'b01 , 2'b01 , 2'b10 , 2'b00 , 2'b00 },
		{ 2'b00 , 2'b00 , 2'b10 , 2'b01 , 2'b01 , 2'b01 , 2'b10 , 2'b10 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b10 , 2'b10 , 2'b01 , 2'b01 , 2'b01 , 2'b10 , 2'b00 , 2'b00 },
		{ 2'b00 , 2'b00 , 2'b10 , 2'b01 , 2'b01 , 2'b01 , 2'b10 , 2'b10 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b10 , 2'b10 , 2'b10 , 2'b01 , 2'b01 , 2'b01 , 2'b10 , 2'b00 , 2'b00 },
		{ 2'b00 , 2'b00 , 2'b10 , 2'b01 , 2'b01 , 2'b01 , 2'b10 , 2'b10 , 2'b10 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b10 , 2'b10 , 2'b10 , 2'b01 , 2'b01 , 2'b01 , 2'b10 , 2'b00 , 2'b00 },
		{ 2'b00 , 2'b00 , 2'b10 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b10 , 2'b10 , 2'b10 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b10 , 2'b10 , 2'b10 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b10 , 2'b00 , 2'b00 },
		{ 2'b00 , 2'b00 , 2'b10 , 2'b10 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b10 , 2'b10 , 2'b10 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b10 , 2'b10 , 2'b10 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b10 , 2'b10 , 2'b00 , 2'b00 },
		{ 2'b00 , 2'b00 , 2'b00 , 2'b10 , 2'b10 , 2'b10 , 2'b10 , 2'b10 , 2'b10 , 2'b10 , 2'b10 , 2'b10 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b10 , 2'b10 , 2'b10 , 2'b10 , 2'b10 , 2'b10 , 2'b10 , 2'b10 , 2'b10 , 2'b00 , 2'b00 , 2'b00 },
		{ 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b10 , 2'b10 , 2'b10 , 2'b10 , 2'b10 , 2'b10 , 2'b10 , 2'b10 , 2'b10 , 2'b10 , 2'b10 , 2'b10 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b10 , 2'b10 , 2'b10 , 2'b10 , 2'b10 , 2'b10 , 2'b10 , 2'b10 , 2'b10 , 2'b10 , 2'b10 , 2'b10 , 2'b00 , 2'b00 , 2'b00 , 2'b00 },
		{ 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b10 , 2'b10 , 2'b10 , 2'b10 , 2'b10 , 2'b11 , 2'b11 , 2'b10 , 2'b10 , 2'b10 , 2'b10 , 2'b10 , 2'b10 , 2'b10 , 2'b10 , 2'b10 , 2'b10 , 2'b11 , 2'b11 , 2'b10 , 2'b10 , 2'b10 , 2'b10 , 2'b10 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 },
		{ 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b10 , 2'b10 , 2'b10 , 2'b10 , 2'b10 , 2'b11 , 2'b11 , 2'b10 , 2'b10 , 2'b10 , 2'b10 , 2'b10 , 2'b10 , 2'b10 , 2'b10 , 2'b10 , 2'b10 , 2'b11 , 2'b11 , 2'b10 , 2'b10 , 2'b10 , 2'b10 , 2'b10 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 },
		{ 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b10 , 2'b10 , 2'b10 , 2'b10 , 2'b11 , 2'b11 , 2'b11 , 2'b10 , 2'b10 , 2'b10 , 2'b10 , 2'b10 , 2'b10 , 2'b10 , 2'b10 , 2'b10 , 2'b10 , 2'b11 , 2'b11 , 2'b11 , 2'b10 , 2'b10 , 2'b10 , 2'b10 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 },
		{ 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b10 , 2'b10 , 2'b11 , 2'b11 , 2'b11 , 2'b11 , 2'b11 , 2'b11 , 2'b11 , 2'b11 , 2'b11 , 2'b11 , 2'b11 , 2'b11 , 2'b11 , 2'b11 , 2'b11 , 2'b11 , 2'b11 , 2'b11 , 2'b10 , 2'b10 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 },
		{ 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b10 , 2'b10 , 2'b11 , 2'b11 , 2'b11 , 2'b11 , 2'b11 , 2'b11 , 2'b10 , 2'b10 , 2'b10 , 2'b10 , 2'b10 , 2'b10 , 2'b11 , 2'b11 , 2'b11 , 2'b11 , 2'b11 , 2'b11 , 2'b10 , 2'b10 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 },
		{ 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b10 , 2'b11 , 2'b11 , 2'b11 , 2'b11 , 2'b11 , 2'b11 , 2'b11 , 2'b11 , 2'b11 , 2'b11 , 2'b11 , 2'b11 , 2'b11 , 2'b11 , 2'b11 , 2'b11 , 2'b11 , 2'b11 , 2'b10 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 },
		{ 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b10 , 2'b10 , 2'b10 , 2'b10 , 2'b10 , 2'b10 , 2'b10 , 2'b10 , 2'b10 , 2'b10 , 2'b10 , 2'b10 , 2'b10 , 2'b10 , 2'b10 , 2'b10 , 2'b10 , 2'b10 , 2'b10 , 2'b10 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 },
		{ 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 },
		{ 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 }
		 },
		{ { 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 },
		{ 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 },
		{ 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b10 , 2'b10 , 2'b10 , 2'b10 , 2'b10 , 2'b10 , 2'b10 , 2'b10 , 2'b10 , 2'b10 , 2'b10 , 2'b10 , 2'b10 , 2'b10 , 2'b10 , 2'b10 , 2'b10 , 2'b10 , 2'b10 , 2'b10 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 },
		{ 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b10 , 2'b11 , 2'b11 , 2'b11 , 2'b11 , 2'b11 , 2'b11 , 2'b11 , 2'b11 , 2'b11 , 2'b11 , 2'b11 , 2'b11 , 2'b11 , 2'b11 , 2'b11 , 2'b11 , 2'b11 , 2'b11 , 2'b10 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 },
		{ 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b10 , 2'b10 , 2'b11 , 2'b11 , 2'b11 , 2'b11 , 2'b11 , 2'b11 , 2'b10 , 2'b10 , 2'b10 , 2'b10 , 2'b10 , 2'b10 , 2'b11 , 2'b11 , 2'b11 , 2'b11 , 2'b11 , 2'b11 , 2'b10 , 2'b10 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 },
		{ 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b10 , 2'b10 , 2'b11 , 2'b11 , 2'b11 , 2'b11 , 2'b11 , 2'b11 , 2'b11 , 2'b11 , 2'b11 , 2'b11 , 2'b11 , 2'b11 , 2'b11 , 2'b11 , 2'b11 , 2'b11 , 2'b11 , 2'b11 , 2'b10 , 2'b10 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 },
		{ 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b10 , 2'b10 , 2'b10 , 2'b10 , 2'b11 , 2'b11 , 2'b11 , 2'b10 , 2'b10 , 2'b10 , 2'b10 , 2'b10 , 2'b10 , 2'b10 , 2'b10 , 2'b10 , 2'b10 , 2'b11 , 2'b11 , 2'b11 , 2'b10 , 2'b10 , 2'b10 , 2'b10 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 },
		{ 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b10 , 2'b10 , 2'b10 , 2'b10 , 2'b10 , 2'b11 , 2'b11 , 2'b10 , 2'b10 , 2'b10 , 2'b10 , 2'b10 , 2'b10 , 2'b10 , 2'b10 , 2'b10 , 2'b10 , 2'b11 , 2'b11 , 2'b10 , 2'b10 , 2'b10 , 2'b10 , 2'b10 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 },
		{ 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b10 , 2'b10 , 2'b10 , 2'b10 , 2'b10 , 2'b11 , 2'b11 , 2'b10 , 2'b10 , 2'b10 , 2'b10 , 2'b10 , 2'b10 , 2'b10 , 2'b10 , 2'b10 , 2'b10 , 2'b11 , 2'b11 , 2'b10 , 2'b10 , 2'b10 , 2'b10 , 2'b10 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 },
		{ 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b10 , 2'b10 , 2'b10 , 2'b10 , 2'b10 , 2'b10 , 2'b10 , 2'b10 , 2'b10 , 2'b10 , 2'b10 , 2'b10 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b10 , 2'b10 , 2'b10 , 2'b10 , 2'b10 , 2'b10 , 2'b10 , 2'b10 , 2'b10 , 2'b10 , 2'b10 , 2'b10 , 2'b00 , 2'b00 , 2'b00 , 2'b00 },
		{ 2'b00 , 2'b00 , 2'b00 , 2'b10 , 2'b10 , 2'b10 , 2'b10 , 2'b10 , 2'b10 , 2'b10 , 2'b10 , 2'b10 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b10 , 2'b10 , 2'b10 , 2'b10 , 2'b10 , 2'b10 , 2'b10 , 2'b10 , 2'b10 , 2'b00 , 2'b00 , 2'b00 },
		{ 2'b00 , 2'b00 , 2'b10 , 2'b10 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b10 , 2'b10 , 2'b10 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b10 , 2'b10 , 2'b10 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b10 , 2'b10 , 2'b00 , 2'b00 },
		{ 2'b00 , 2'b00 , 2'b10 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b10 , 2'b10 , 2'b10 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b10 , 2'b10 , 2'b10 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b10 , 2'b00 , 2'b00 },
		{ 2'b00 , 2'b00 , 2'b10 , 2'b01 , 2'b01 , 2'b01 , 2'b10 , 2'b10 , 2'b10 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b10 , 2'b10 , 2'b10 , 2'b01 , 2'b01 , 2'b01 , 2'b10 , 2'b00 , 2'b00 },
		{ 2'b00 , 2'b00 , 2'b10 , 2'b01 , 2'b01 , 2'b01 , 2'b10 , 2'b10 , 2'b10 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b10 , 2'b10 , 2'b01 , 2'b01 , 2'b01 , 2'b10 , 2'b00 , 2'b00 },
		{ 2'b00 , 2'b00 , 2'b10 , 2'b01 , 2'b01 , 2'b01 , 2'b10 , 2'b10 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b10 , 2'b10 , 2'b01 , 2'b01 , 2'b01 , 2'b10 , 2'b00 , 2'b00 },
		{ 2'b00 , 2'b00 , 2'b10 , 2'b01 , 2'b01 , 2'b01 , 2'b10 , 2'b10 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b10 , 2'b10 , 2'b01 , 2'b01 , 2'b01 , 2'b10 , 2'b00 , 2'b00 },
		{ 2'b00 , 2'b00 , 2'b10 , 2'b01 , 2'b01 , 2'b01 , 2'b10 , 2'b10 , 2'b10 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b10 , 2'b10 , 2'b01 , 2'b01 , 2'b01 , 2'b10 , 2'b00 , 2'b00 },
		{ 2'b00 , 2'b00 , 2'b10 , 2'b01 , 2'b01 , 2'b01 , 2'b10 , 2'b10 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b10 , 2'b10 , 2'b01 , 2'b01 , 2'b01 , 2'b10 , 2'b00 , 2'b00 },
		{ 2'b00 , 2'b00 , 2'b10 , 2'b01 , 2'b01 , 2'b01 , 2'b10 , 2'b10 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b10 , 2'b10 , 2'b01 , 2'b01 , 2'b10 , 2'b10 , 2'b00 , 2'b00 },
		{ 2'b00 , 2'b00 , 2'b10 , 2'b01 , 2'b01 , 2'b01 , 2'b10 , 2'b10 , 2'b10 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b10 , 2'b10 , 2'b10 , 2'b01 , 2'b10 , 2'b10 , 2'b10 , 2'b00 , 2'b00 },
		{ 2'b00 , 2'b00 , 2'b10 , 2'b01 , 2'b01 , 2'b01 , 2'b10 , 2'b10 , 2'b10 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b10 , 2'b10 , 2'b10 , 2'b10 , 2'b10 , 2'b00 , 2'b00 , 2'b00 , 2'b00 },
		{ 2'b00 , 2'b00 , 2'b10 , 2'b01 , 2'b01 , 2'b01 , 2'b10 , 2'b10 , 2'b10 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b10 , 2'b10 , 2'b10 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 },
		{ 2'b00 , 2'b00 , 2'b10 , 2'b01 , 2'b01 , 2'b01 , 2'b10 , 2'b10 , 2'b10 , 2'b10 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b10 , 2'b10 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 },
		{ 2'b10 , 2'b10 , 2'b10 , 2'b01 , 2'b01 , 2'b01 , 2'b10 , 2'b10 , 2'b11 , 2'b10 , 2'b10 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b10 , 2'b10 , 2'b10 , 2'b10 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 },
		{ 2'b10 , 2'b11 , 2'b10 , 2'b10 , 2'b01 , 2'b01 , 2'b10 , 2'b10 , 2'b11 , 2'b11 , 2'b10 , 2'b10 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b10 , 2'b10 , 2'b10 , 2'b11 , 2'b10 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 },
		{ 2'b10 , 2'b11 , 2'b11 , 2'b10 , 2'b01 , 2'b01 , 2'b01 , 2'b10 , 2'b11 , 2'b11 , 2'b10 , 2'b10 , 2'b10 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b10 , 2'b10 , 2'b10 , 2'b11 , 2'b11 , 2'b10 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 },
		{ 2'b10 , 2'b11 , 2'b11 , 2'b10 , 2'b10 , 2'b01 , 2'b01 , 2'b10 , 2'b11 , 2'b11 , 2'b10 , 2'b00 , 2'b10 , 2'b10 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b10 , 2'b10 , 2'b11 , 2'b11 , 2'b11 , 2'b11 , 2'b10 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 },
		{ 2'b10 , 2'b10 , 2'b10 , 2'b10 , 2'b10 , 2'b10 , 2'b01 , 2'b10 , 2'b11 , 2'b11 , 2'b10 , 2'b00 , 2'b10 , 2'b10 , 2'b10 , 2'b10 , 2'b10 , 2'b10 , 2'b10 , 2'b10 , 2'b10 , 2'b10 , 2'b10 , 2'b10 , 2'b10 , 2'b10 , 2'b10 , 2'b10 , 2'b11 , 2'b11 , 2'b11 , 2'b11 , 2'b10 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 },
		{ 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b10 , 2'b01 , 2'b10 , 2'b11 , 2'b11 , 2'b10 , 2'b00 , 2'b00 , 2'b10 , 2'b10 , 2'b10 , 2'b10 , 2'b10 , 2'b10 , 2'b10 , 2'b10 , 2'b10 , 2'b10 , 2'b10 , 2'b10 , 2'b10 , 2'b11 , 2'b11 , 2'b11 , 2'b11 , 2'b11 , 2'b11 , 2'b10 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 },
		{ 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b10 , 2'b10 , 2'b10 , 2'b11 , 2'b11 , 2'b10 , 2'b00 , 2'b00 , 2'b10 , 2'b11 , 2'b11 , 2'b11 , 2'b11 , 2'b11 , 2'b11 , 2'b11 , 2'b10 , 2'b00 , 2'b10 , 2'b10 , 2'b11 , 2'b11 , 2'b11 , 2'b11 , 2'b11 , 2'b11 , 2'b10 , 2'b10 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 },
		{ 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b10 , 2'b10 , 2'b11 , 2'b11 , 2'b10 , 2'b00 , 2'b00 , 2'b10 , 2'b10 , 2'b11 , 2'b11 , 2'b11 , 2'b11 , 2'b11 , 2'b11 , 2'b10 , 2'b00 , 2'b00 , 2'b10 , 2'b10 , 2'b11 , 2'b11 , 2'b11 , 2'b11 , 2'b10 , 2'b10 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 },
		{ 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b10 , 2'b11 , 2'b11 , 2'b10 , 2'b00 , 2'b00 , 2'b00 , 2'b10 , 2'b10 , 2'b11 , 2'b11 , 2'b11 , 2'b11 , 2'b10 , 2'b10 , 2'b00 , 2'b00 , 2'b00 , 2'b10 , 2'b10 , 2'b10 , 2'b10 , 2'b10 , 2'b10 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 },
		{ 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b10 , 2'b11 , 2'b11 , 2'b10 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b10 , 2'b10 , 2'b10 , 2'b10 , 2'b10 , 2'b10 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 },
		{ 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b10 , 2'b11 , 2'b11 , 2'b10 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 },
		{ 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b10 , 2'b11 , 2'b11 , 2'b10 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 },
		{ 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b10 , 2'b11 , 2'b11 , 2'b10 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 },
		{ 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b10 , 2'b11 , 2'b11 , 2'b10 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 },
		{ 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b10 , 2'b10 , 2'b11 , 2'b11 , 2'b10 , 2'b10 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 },
		{ 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b10 , 2'b10 , 2'b10 , 2'b10 , 2'b10 , 2'b10 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 }
		 },
		{ { 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b10 , 2'b10 , 2'b10 , 2'b10 , 2'b10 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 },
		{ 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b10 , 2'b11 , 2'b11 , 2'b11 , 2'b10 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 },
		{ 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b10 , 2'b11 , 2'b11 , 2'b10 , 2'b10 , 2'b10 , 2'b10 , 2'b10 , 2'b10 , 2'b10 , 2'b10 , 2'b10 , 2'b10 , 2'b10 , 2'b10 , 2'b10 , 2'b10 , 2'b10 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 },
		{ 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b10 , 2'b10 , 2'b10 , 2'b10 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b10 , 2'b10 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 },
		{ 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b10 , 2'b10 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b10 , 2'b10 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 },
		{ 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b10 , 2'b10 , 2'b10 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b10 , 2'b10 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 },
		{ 2'b10 , 2'b10 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b10 , 2'b10 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b10 , 2'b10 , 2'b10 , 2'b10 , 2'b10 , 2'b10 , 2'b10 , 2'b10 , 2'b10 , 2'b10 , 2'b10 , 2'b10 , 2'b10 , 2'b01 , 2'b01 , 2'b10 , 2'b10 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 },
		{ 2'b10 , 2'b10 , 2'b10 , 2'b10 , 2'b10 , 2'b10 , 2'b10 , 2'b10 , 2'b10 , 2'b10 , 2'b10 , 2'b10 , 2'b10 , 2'b10 , 2'b10 , 2'b10 , 2'b10 , 2'b10 , 2'b10 , 2'b10 , 2'b10 , 2'b10 , 2'b10 , 2'b10 , 2'b10 , 2'b10 , 2'b10 , 2'b10 , 2'b01 , 2'b10 , 2'b10 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 },
		{ 2'b10 , 2'b11 , 2'b11 , 2'b11 , 2'b11 , 2'b11 , 2'b11 , 2'b11 , 2'b11 , 2'b11 , 2'b11 , 2'b11 , 2'b11 , 2'b11 , 2'b11 , 2'b11 , 2'b10 , 2'b10 , 2'b10 , 2'b10 , 2'b01 , 2'b01 , 2'b10 , 2'b01 , 2'b01 , 2'b10 , 2'b10 , 2'b10 , 2'b10 , 2'b10 , 2'b10 , 2'b10 , 2'b10 , 2'b10 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 },
		{ 2'b10 , 2'b11 , 2'b11 , 2'b11 , 2'b11 , 2'b11 , 2'b11 , 2'b11 , 2'b11 , 2'b11 , 2'b11 , 2'b11 , 2'b11 , 2'b11 , 2'b11 , 2'b10 , 2'b10 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b10 , 2'b10 , 2'b10 , 2'b10 , 2'b10 , 2'b10 , 2'b10 , 2'b10 , 2'b10 , 2'b00 , 2'b00 , 2'b00 , 2'b00 },
		{ 2'b10 , 2'b10 , 2'b10 , 2'b10 , 2'b10 , 2'b10 , 2'b10 , 2'b10 , 2'b10 , 2'b10 , 2'b10 , 2'b10 , 2'b10 , 2'b10 , 2'b10 , 2'b10 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b10 , 2'b10 , 2'b10 , 2'b10 , 2'b10 , 2'b10 , 2'b10 , 2'b10 , 2'b10 , 2'b10 , 2'b00 , 2'b00 },
		{ 2'b10 , 2'b10 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b10 , 2'b10 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b10 , 2'b10 , 2'b10 , 2'b10 , 2'b10 , 2'b11 , 2'b11 , 2'b11 , 2'b10 , 2'b00 , 2'b00 },
		{ 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b10 , 2'b10 , 2'b10 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b10 , 2'b10 , 2'b10 , 2'b11 , 2'b11 , 2'b11 , 2'b11 , 2'b10 , 2'b00 , 2'b00 },
		{ 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b10 , 2'b10 , 2'b10 , 2'b10 , 2'b10 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b10 , 2'b11 , 2'b11 , 2'b11 , 2'b11 , 2'b11 , 2'b11 , 2'b10 , 2'b00 , 2'b00 },
		{ 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b10 , 2'b10 , 2'b11 , 2'b10 , 2'b10 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b10 , 2'b11 , 2'b11 , 2'b11 , 2'b11 , 2'b11 , 2'b11 , 2'b10 , 2'b00 , 2'b00 },
		{ 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b10 , 2'b10 , 2'b11 , 2'b11 , 2'b10 , 2'b10 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b10 , 2'b10 , 2'b10 , 2'b10 , 2'b11 , 2'b11 , 2'b11 , 2'b10 , 2'b00 , 2'b00 },
		{ 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b10 , 2'b11 , 2'b11 , 2'b11 , 2'b10 , 2'b10 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b10 , 2'b10 , 2'b10 , 2'b11 , 2'b11 , 2'b11 , 2'b10 , 2'b00 , 2'b00 },
		{ 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b10 , 2'b11 , 2'b11 , 2'b11 , 2'b10 , 2'b10 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b10 , 2'b10 , 2'b10 , 2'b11 , 2'b10 , 2'b11 , 2'b10 , 2'b00 , 2'b00 },
		{ 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b10 , 2'b11 , 2'b11 , 2'b11 , 2'b10 , 2'b10 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b10 , 2'b10 , 2'b10 , 2'b11 , 2'b10 , 2'b11 , 2'b10 , 2'b00 , 2'b00 },
		{ 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b10 , 2'b11 , 2'b11 , 2'b11 , 2'b10 , 2'b10 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b10 , 2'b10 , 2'b10 , 2'b11 , 2'b10 , 2'b11 , 2'b10 , 2'b00 , 2'b00 },
		{ 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 ,  2'b10 , 2'b10 , 2'b11 , 2'b11 , 2'b10 , 2'b10 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b10 , 2'b10 , 2'b10 , 2'b11 , 2'b10 , 2'b11 , 2'b10 , 2'b00 , 2'b00 },
		{ 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b10 , 2'b10 , 2'b10 , 2'b10 , 2'b10 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b10 , 2'b10 , 2'b10 , 2'b11 , 2'b10 , 2'b11 , 2'b10 , 2'b00 , 2'b00 },
		{ 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b10 , 2'b10 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b10 , 2'b10 , 2'b10 , 2'b11 , 2'b10 , 2'b11 , 2'b10 , 2'b00 , 2'b00 },
		{ 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b10 , 2'b10 , 2'b10 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b10 , 2'b10 , 2'b10 , 2'b11 , 2'b11 , 2'b11 , 2'b10 , 2'b00 , 2'b00 },
		{ 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b10 , 2'b10 , 2'b10 , 2'b10 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b10 , 2'b10 , 2'b10 , 2'b10 , 2'b11 , 2'b11 , 2'b11 , 2'b10 , 2'b00 , 2'b00 },
		{ 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b10 , 2'b10 , 2'b11 , 2'b10 , 2'b10 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b10 , 2'b11 , 2'b11 , 2'b11 , 2'b11 , 2'b11 , 2'b11 , 2'b10 , 2'b00 , 2'b00 },
		{ 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b10 , 2'b11 , 2'b11 , 2'b11 , 2'b10 , 2'b10 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b10 , 2'b11 , 2'b11 , 2'b11 , 2'b11 , 2'b11 , 2'b11 , 2'b10 , 2'b00 , 2'b00 },
		{ 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b10 , 2'b11 , 2'b11 , 2'b11 , 2'b10 , 2'b10 , 2'b10 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b10 , 2'b10 , 2'b10 , 2'b11 , 2'b11 , 2'b11 , 2'b11 , 2'b10 , 2'b00 , 2'b00 },
		{ 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b10 , 2'b11 , 2'b11 , 2'b11 , 2'b11 , 2'b11 , 2'b10 , 2'b10 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b10 , 2'b10 , 2'b10 , 2'b10 , 2'b10 , 2'b11 , 2'b11 , 2'b11 , 2'b10 , 2'b00 , 2'b00 },
		{ 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b10 , 2'b11 , 2'b11 , 2'b11 , 2'b11 , 2'b11 , 2'b10 , 2'b10 , 2'b10 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b10 , 2'b10 , 2'b10 , 2'b10 , 2'b10 , 2'b10 , 2'b10 , 2'b10 , 2'b10 , 2'b10 , 2'b00 , 2'b00 },
		{ 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b10 , 2'b10 , 2'b11 , 2'b11 , 2'b11 , 2'b11 , 2'b11 , 2'b10 , 2'b10 , 2'b10 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b10 , 2'b10 , 2'b10 , 2'b10 , 2'b10 , 2'b10 , 2'b10 , 2'b10 , 2'b10 , 2'b00 , 2'b00 , 2'b00 , 2'b00 },
		{ 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b10 , 2'b10 , 2'b11 , 2'b11 , 2'b11 , 2'b11 , 2'b11 , 2'b10 , 2'b10 , 2'b10 , 2'b10 , 2'b10 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b10 , 2'b10 , 2'b10 , 2'b10 , 2'b10 , 2'b10 , 2'b10 , 2'b10 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 },
		{ 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b10 , 2'b10 , 2'b10 , 2'b10 , 2'b10 , 2'b10 , 2'b10 , 2'b00 , 2'b10 , 2'b10 , 2'b10 , 2'b10 , 2'b10 , 2'b10 , 2'b10 , 2'b10 , 2'b10 , 2'b10 , 2'b10 , 2'b01 , 2'b10 , 2'b10 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 },
		{ 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b10 , 2'b10 , 2'b10 , 2'b10 , 2'b10 , 2'b10 , 2'b10 , 2'b10 , 2'b10 , 2'b10 , 2'b01 , 2'b01 , 2'b10 , 2'b10 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 },
		{ 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b10 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b10 , 2'b10 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 },
		{ 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b10 , 2'b10 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b10 , 2'b10 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 },
		{ 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b10 , 2'b10 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b10 , 2'b10 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 },
		{ 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b10 , 2'b10 , 2'b10 , 2'b10 , 2'b10 , 2'b10 , 2'b10 , 2'b10 , 2'b10 , 2'b10 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 },
		{ 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 },
		{ 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 }
		 },
		{ { 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 },
		{ 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 },
		{ 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b10 , 2'b10 , 2'b10 , 2'b10 , 2'b10 , 2'b10 , 2'b10 , 2'b10 , 2'b10 , 2'b10 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 },
		{ 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b10 , 2'b10 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b10 , 2'b10 , 2'b01 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 },
		{ 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b10 , 2'b10 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b10 , 2'b10 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 },
		{ 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b10 , 2'b10 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b10 , 2'b01 , 2'b10 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 },
		{ 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b10 , 2'b10 , 2'b01 , 2'b01 , 2'b10 , 2'b10 , 2'b10 , 2'b10 , 2'b10 , 2'b10 , 2'b10 , 2'b10 , 2'b10 , 2'b10 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 },
		{ 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b10 , 2'b10 , 2'b01 , 2'b10 , 2'b10 , 2'b10 , 2'b10 , 2'b10 , 2'b10 , 2'b10 , 2'b10 , 2'b10 , 2'b10 , 2'b10 , 2'b00 , 2'b10 , 2'b10 , 2'b10 , 2'b10 , 2'b10 , 2'b10 , 2'b10 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 },
		{ 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b10 , 2'b10 , 2'b10 , 2'b10 , 2'b10 , 2'b10 , 2'b10 , 2'b10 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b10 , 2'b10 , 2'b10 , 2'b10 , 2'b10 , 2'b11 , 2'b11 , 2'b11 , 2'b11 , 2'b11 , 2'b10 , 2'b10 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 },
		{ 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b10 , 2'b10 , 2'b10 , 2'b10 , 2'b10 , 2'b10 , 2'b10 , 2'b10 , 2'b10 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b10 , 2'b10 , 2'b10 , 2'b11 , 2'b11 , 2'b11 , 2'b11 , 2'b11 , 2'b10 , 2'b10 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 },
		{ 2'b00 , 2'b00 , 2'b10 , 2'b10 , 2'b10 , 2'b10 , 2'b10 , 2'b10 , 2'b10 , 2'b10 , 2'b10 , 2'b10 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b10 , 2'b10 , 2'b10 , 2'b11 , 2'b11 , 2'b11 , 2'b11 , 2'b11 , 2'b10 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 },
		{ 2'b00 , 2'b00 , 2'b10 , 2'b11 , 2'b11 , 2'b11 , 2'b10 , 2'b10 , 2'b10 , 2'b10 , 2'b10 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b10 , 2'b10 , 2'b11 , 2'b11 , 2'b11 , 2'b11 , 2'b11 , 2'b10 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 },
		{ 2'b00 , 2'b00 , 2'b10 , 2'b11 , 2'b11 , 2'b11 , 2'b11 , 2'b10 , 2'b10 , 2'b10 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b10 , 2'b10 , 2'b10 , 2'b11 , 2'b11 , 2'b11 , 2'b10 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 },
		{ 2'b00 , 2'b00 , 2'b10 , 2'b11 , 2'b11 , 2'b11 , 2'b11 , 2'b11 , 2'b11 , 2'b10 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b10 , 2'b10 , 2'b11 , 2'b11 , 2'b11 , 2'b10 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 },
		{ 2'b00 , 2'b00 , 2'b10 , 2'b11 , 2'b11 , 2'b11 , 2'b11 , 2'b11 , 2'b11 , 2'b10 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b10 , 2'b10 , 2'b11 , 2'b10 , 2'b10 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 },
		{ 2'b00 , 2'b00 , 2'b10 , 2'b11 , 2'b11 , 2'b11 , 2'b10 , 2'b10 , 2'b10 , 2'b10 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b10 , 2'b10 , 2'b10 , 2'b10 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 },
		{ 2'b00 , 2'b00 , 2'b10 , 2'b11 , 2'b11 , 2'b11 , 2'b10 , 2'b10 , 2'b10 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b10 , 2'b10 , 2'b10 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 },
		{ 2'b00 , 2'b00 , 2'b10 , 2'b11 , 2'b10 , 2'b11 , 2'b10 , 2'b10 , 2'b10 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b10 , 2'b10 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 },
		{ 2'b00 , 2'b00 , 2'b10 , 2'b11 , 2'b10 , 2'b11 , 2'b10 , 2'b10 , 2'b10 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b10 , 2'b10 , 2'b10 , 2'b10 , 2'b10 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 },
		{ 2'b00 , 2'b00 , 2'b10 , 2'b11 , 2'b10 , 2'b11 , 2'b10 , 2'b10 , 2'b10 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b10 , 2'b10 , 2'b11 , 2'b11 , 2'b10 , 2'b10 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 },
		{ 2'b00 , 2'b00 , 2'b10 , 2'b11 , 2'b10 , 2'b11 , 2'b10 , 2'b10 , 2'b10 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b10 , 2'b10 , 2'b11 , 2'b11 , 2'b11 , 2'b10 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 },
		{ 2'b00 , 2'b00 , 2'b10 , 2'b11 , 2'b10 , 2'b11 , 2'b10 , 2'b10 , 2'b10 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b10 , 2'b10 , 2'b11 , 2'b11 , 2'b11 , 2'b10 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 },
		{ 2'b00 , 2'b00 , 2'b10 , 2'b11 , 2'b10 , 2'b11 , 2'b10 , 2'b10 , 2'b10 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b10 , 2'b10 , 2'b11 , 2'b11 , 2'b11 , 2'b10 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 },
		{ 2'b00 , 2'b00 , 2'b10 , 2'b11 , 2'b11 , 2'b11 , 2'b10 , 2'b10 , 2'b10 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b10 , 2'b10 , 2'b11 , 2'b11 , 2'b11 , 2'b10 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 },
		{ 2'b00 , 2'b00 , 2'b10 , 2'b11 , 2'b11 , 2'b11 , 2'b10 , 2'b10 , 2'b10 , 2'b10 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b10 , 2'b10 , 2'b11 , 2'b11 , 2'b10 , 2'b10 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 },
		{ 2'b00 , 2'b00 , 2'b10 , 2'b11 , 2'b11 , 2'b11 , 2'b11 , 2'b11 , 2'b11 , 2'b10 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b10 , 2'b10 , 2'b11 , 2'b10 , 2'b10 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 },
		{ 2'b00 , 2'b00 , 2'b10 , 2'b11 , 2'b11 , 2'b11 , 2'b11 , 2'b11 , 2'b11 , 2'b10 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b10 , 2'b10 , 2'b10 , 2'b10 , 2'b10 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 },
		{ 2'b00 , 2'b00 , 2'b10 , 2'b11 , 2'b11 , 2'b11 , 2'b11 , 2'b10 , 2'b10 , 2'b10 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b10 , 2'b10 , 2'b10 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 },
		{ 2'b00 , 2'b00 , 2'b10 , 2'b11 , 2'b11 , 2'b11 , 2'b10 , 2'b10 , 2'b10 , 2'b10 , 2'b10 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b10 , 2'b10 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b10 , 2'b10 },
		{ 2'b00 , 2'b00 , 2'b10 , 2'b10 , 2'b10 , 2'b10 , 2'b10 , 2'b10 , 2'b10 , 2'b10 , 2'b10 , 2'b10 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b10 , 2'b10 , 2'b10 , 2'b10 , 2'b10 , 2'b10 , 2'b10 , 2'b10 , 2'b10 , 2'b10 , 2'b10 , 2'b10 , 2'b10 , 2'b10 , 2'b10 , 2'b10 },
		{ 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b10 , 2'b10 , 2'b10 , 2'b10 , 2'b10 , 2'b10 , 2'b10 , 2'b10 , 2'b10 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b10 , 2'b10 , 2'b11 , 2'b11 , 2'b11 , 2'b11 , 2'b11 , 2'b11 , 2'b11 , 2'b11 , 2'b11 , 2'b11 , 2'b11 , 2'b11 , 2'b11 , 2'b11 , 2'b10 },
		{ 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b10 , 2'b10 , 2'b10 , 2'b10 , 2'b10 , 2'b10 , 2'b10 , 2'b10 , 2'b10 , 2'b01 , 2'b01 , 2'b10 , 2'b01 , 2'b01 , 2'b10 , 2'b10 , 2'b10 , 2'b10 , 2'b11 , 2'b11 , 2'b11 , 2'b11 , 2'b11 , 2'b11 , 2'b11 , 2'b11 , 2'b11 , 2'b11 , 2'b11 , 2'b11 , 2'b11 , 2'b11 , 2'b11 , 2'b10 },
		{ 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b10 , 2'b10 , 2'b01 , 2'b10 , 2'b10 , 2'b10 , 2'b10 , 2'b10 , 2'b10 , 2'b10 , 2'b10 , 2'b10 , 2'b10 , 2'b10 , 2'b10 , 2'b10 , 2'b10 , 2'b10 , 2'b10 , 2'b10 , 2'b10 , 2'b10 , 2'b10 , 2'b10 , 2'b10 , 2'b10 , 2'b10 , 2'b10 , 2'b10 , 2'b10 , 2'b10 },
		{ 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b10 , 2'b10 , 2'b01 , 2'b01 , 2'b10 , 2'b10 , 2'b10 , 2'b10 , 2'b10 , 2'b10 , 2'b10 , 2'b10 , 2'b10 , 2'b10 , 2'b10 , 2'b10 , 2'b10 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b10 , 2'b10 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 },
		{ 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b10 , 2'b10 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b10 , 2'b10 , 2'b10 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 },
		{ 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b01 , 2'b01 , 2'b10 , 2'b10 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b10 , 2'b10 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 },
		{ 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b10 , 2'b10 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b01 , 2'b10 , 2'b10 , 2'b10 , 2'b10 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 },
		{ 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b10 , 2'b10 , 2'b10 , 2'b10 , 2'b10 , 2'b10 , 2'b10 , 2'b10 , 2'b10 , 2'b10 , 2'b10 , 2'b10 , 2'b10 , 2'b10 , 2'b10 , 2'b11 , 2'b11 , 2'b10 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 },
		{ 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b10 , 2'b11 , 2'b11 , 2'b11 , 2'b10 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 },
		{ 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b10 , 2'b10 , 2'b10 , 2'b10 , 2'b10 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 , 2'b00 }}};

    assign data = en ? rom[dir][y][x] : 2'b00;

endmodule