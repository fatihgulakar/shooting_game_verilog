//----------------------------------------------------------------------------------
//-- Object file that contains pixel data of player characters
//----------------------------------------------------------------------------------


module obj_p(
    input [5:0]  x,
    input [5:0]  y,
    input [1:0]  dir, //0 up, 1 down, 2 left ,3 right
    input        en,
    output [1:0] data
);
 
reg [0:1] rom [1:0][0:39][0:39];
//	type arr is array ( 0 to 3 , 0 to 39 , 0 to 39 ) of std_logic_vector( 1 downto 0 );
initial begin
 rom[0][0][0] = 2'b00;	 rom[0][1][0] = 2'b00;	 rom[0][2][0] = 2'b00;	 rom[0][3][0] = 2'b00;	 rom[0][4][0] = 2'b00;	 rom[0][5][0] = 2'b00;	 rom[0][6][0] = 2'b00;	 rom[0][7][0] = 2'b00;	 rom[0][8][0] = 2'b00;	 rom[0][9][0] = 2'b00;	 rom[0][10][0] = 2'b00;	 rom[0][11][0] = 2'b00;	 rom[0][12][0] = 2'b00;	 rom[0][13][0] = 2'b00;	 rom[0][14][0] = 2'b00;	 rom[0][15][0] = 2'b00;	 rom[0][16][0] = 2'b00;	 rom[0][17][0] = 2'b00;	 rom[0][18][0] = 2'b00;	 rom[0][19][0] = 2'b00;	 rom[0][20][0] = 2'b00;	 rom[0][21][0] = 2'b00;	 rom[0][22][0] = 2'b00;	 rom[0][23][0] = 2'b00;	 rom[0][24][0] = 2'b00;	 rom[0][25][0] = 2'b00;	 rom[0][26][0] = 2'b00;	 rom[0][27][0] = 2'b00;	 rom[0][28][0] = 2'b10;	 rom[0][29][0] = 2'b10;	 rom[0][30][0] = 2'b10;	 rom[0][31][0] = 2'b10;	 rom[0][32][0] = 2'b10;	 rom[0][33][0] = 2'b10;	 rom[0][34][0] = 2'b00;	 rom[0][35][0] = 2'b00;	 rom[0][36][0] = 2'b00;	 rom[0][37][0] = 2'b00;	 rom[0][38][0] = 2'b00;	 rom[0][39][0] = 2'b00;
 rom[0][0][1] = 2'b00;	 rom[0][1][1] = 2'b00;	 rom[0][2][1] = 2'b00;	 rom[0][3][1] = 2'b00;	 rom[0][4][1] = 2'b00;	 rom[0][5][1] = 2'b00;	 rom[0][6][1] = 2'b00;	 rom[0][7][1] = 2'b00;	 rom[0][8][1] = 2'b00;	 rom[0][9][1] = 2'b00;	 rom[0][10][1] = 2'b00;	 rom[0][11][1] = 2'b00;	 rom[0][12][1] = 2'b00;	 rom[0][13][1] = 2'b00;	 rom[0][14][1] = 2'b00;	 rom[0][15][1] = 2'b00;	 rom[0][16][1] = 2'b00;	 rom[0][17][1] = 2'b00;	 rom[0][18][1] = 2'b00;	 rom[0][19][1] = 2'b00;	 rom[0][20][1] = 2'b00;	 rom[0][21][1] = 2'b00;	 rom[0][22][1] = 2'b00;	 rom[0][23][1] = 2'b00;	 rom[0][24][1] = 2'b00;	 rom[0][25][1] = 2'b00;	 rom[0][26][1] = 2'b00;	 rom[0][27][1] = 2'b00;	 rom[0][28][1] = 2'b10;	 rom[0][29][1] = 2'b10;	 rom[0][30][1] = 2'b11;	 rom[0][31][1] = 2'b11;	 rom[0][32][1] = 2'b10;	 rom[0][33][1] = 2'b10;	 rom[0][34][1] = 2'b00;	 rom[0][35][1] = 2'b00;	 rom[0][36][1] = 2'b00;	 rom[0][37][1] = 2'b00;	 rom[0][38][1] = 2'b00;	 rom[0][39][1] = 2'b00;
 rom[0][0][2] = 2'b00;	 rom[0][1][2] = 2'b00;	 rom[0][2][2] = 2'b00;	 rom[0][3][2] = 2'b00;	 rom[0][4][2] = 2'b00;	 rom[0][5][2] = 2'b00;	 rom[0][6][2] = 2'b00;	 rom[0][7][2] = 2'b00;	 rom[0][8][2] = 2'b00;	 rom[0][9][2] = 2'b00;	 rom[0][10][2] = 2'b00;	 rom[0][11][2] = 2'b00;	 rom[0][12][2] = 2'b00;	 rom[0][13][2] = 2'b00;	 rom[0][14][2] = 2'b00;	 rom[0][15][2] = 2'b00;	 rom[0][16][2] = 2'b00;	 rom[0][17][2] = 2'b00;	 rom[0][18][2] = 2'b00;	 rom[0][19][2] = 2'b00;	 rom[0][20][2] = 2'b00;	 rom[0][21][2] = 2'b00;	 rom[0][22][2] = 2'b00;	 rom[0][23][2] = 2'b00;	 rom[0][24][2] = 2'b00;	 rom[0][25][2] = 2'b00;	 rom[0][26][2] = 2'b00;	 rom[0][27][2] = 2'b00;	 rom[0][28][2] = 2'b00;	 rom[0][29][2] = 2'b10;	 rom[0][30][2] = 2'b11;	 rom[0][31][2] = 2'b11;	 rom[0][32][2] = 2'b10;	 rom[0][33][2] = 2'b00;	 rom[0][34][2] = 2'b00;	 rom[0][35][2] = 2'b00;	 rom[0][36][2] = 2'b00;	 rom[0][37][2] = 2'b00;	 rom[0][38][2] = 2'b00;	 rom[0][39][2] = 2'b00;
 rom[0][0][3] = 2'b00;	 rom[0][1][3] = 2'b00;	 rom[0][2][3] = 2'b00;	 rom[0][3][3] = 2'b00;	 rom[0][4][3] = 2'b00;	 rom[0][5][3] = 2'b00;	 rom[0][6][3] = 2'b00;	 rom[0][7][3] = 2'b00;	 rom[0][8][3] = 2'b00;	 rom[0][9][3] = 2'b00;	 rom[0][10][3] = 2'b00;	 rom[0][11][3] = 2'b00;	 rom[0][12][3] = 2'b00;	 rom[0][13][3] = 2'b00;	 rom[0][14][3] = 2'b00;	 rom[0][15][3] = 2'b00;	 rom[0][16][3] = 2'b00;	 rom[0][17][3] = 2'b00;	 rom[0][18][3] = 2'b00;	 rom[0][19][3] = 2'b00;	 rom[0][20][3] = 2'b00;	 rom[0][21][3] = 2'b00;	 rom[0][22][3] = 2'b00;	 rom[0][23][3] = 2'b00;	 rom[0][24][3] = 2'b00;	 rom[0][25][3] = 2'b00;	 rom[0][26][3] = 2'b00;	 rom[0][27][3] = 2'b00;	 rom[0][28][3] = 2'b00;	 rom[0][29][3] = 2'b10;	 rom[0][30][3] = 2'b11;	 rom[0][31][3] = 2'b11;	 rom[0][32][3] = 2'b10;	 rom[0][33][3] = 2'b00;	 rom[0][34][3] = 2'b00;	 rom[0][35][3] = 2'b00;	 rom[0][36][3] = 2'b00;	 rom[0][37][3] = 2'b00;	 rom[0][38][3] = 2'b00;	 rom[0][39][3] = 2'b00;
 rom[0][0][4] = 2'b00;	 rom[0][1][4] = 2'b00;	 rom[0][2][4] = 2'b00;	 rom[0][3][4] = 2'b00;	 rom[0][4][4] = 2'b00;	 rom[0][5][4] = 2'b00;	 rom[0][6][4] = 2'b00;	 rom[0][7][4] = 2'b00;	 rom[0][8][4] = 2'b00;	 rom[0][9][4] = 2'b00;	 rom[0][10][4] = 2'b00;	 rom[0][11][4] = 2'b00;	 rom[0][12][4] = 2'b00;	 rom[0][13][4] = 2'b00;	 rom[0][14][4] = 2'b00;	 rom[0][15][4] = 2'b00;	 rom[0][16][4] = 2'b00;	 rom[0][17][4] = 2'b00;	 rom[0][18][4] = 2'b00;	 rom[0][19][4] = 2'b00;	 rom[0][20][4] = 2'b00;	 rom[0][21][4] = 2'b00;	 rom[0][22][4] = 2'b00;	 rom[0][23][4] = 2'b00;	 rom[0][24][4] = 2'b00;	 rom[0][25][4] = 2'b00;	 rom[0][26][4] = 2'b00;	 rom[0][27][4] = 2'b00;	 rom[0][28][4] = 2'b00;	 rom[0][29][4] = 2'b10;	 rom[0][30][4] = 2'b11;	 rom[0][31][4] = 2'b11;	 rom[0][32][4] = 2'b10;	 rom[0][33][4] = 2'b00;	 rom[0][34][4] = 2'b00;	 rom[0][35][4] = 2'b00;	 rom[0][36][4] = 2'b00;	 rom[0][37][4] = 2'b00;	 rom[0][38][4] = 2'b00;	 rom[0][39][4] = 2'b00;
 rom[0][0][5] = 2'b00;	 rom[0][1][5] = 2'b00;	 rom[0][2][5] = 2'b00;	 rom[0][3][5] = 2'b00;	 rom[0][4][5] = 2'b00;	 rom[0][5][5] = 2'b00;	 rom[0][6][5] = 2'b00;	 rom[0][7][5] = 2'b00;	 rom[0][8][5] = 2'b00;	 rom[0][9][5] = 2'b00;	 rom[0][10][5] = 2'b00;	 rom[0][11][5] = 2'b00;	 rom[0][12][5] = 2'b00;	 rom[0][13][5] = 2'b00;	 rom[0][14][5] = 2'b00;	 rom[0][15][5] = 2'b00;	 rom[0][16][5] = 2'b00;	 rom[0][17][5] = 2'b00;	 rom[0][18][5] = 2'b00;	 rom[0][19][5] = 2'b00;	 rom[0][20][5] = 2'b00;	 rom[0][21][5] = 2'b00;	 rom[0][22][5] = 2'b00;	 rom[0][23][5] = 2'b00;	 rom[0][24][5] = 2'b00;	 rom[0][25][5] = 2'b00;	 rom[0][26][5] = 2'b00;	 rom[0][27][5] = 2'b00;	 rom[0][28][5] = 2'b00;	 rom[0][29][5] = 2'b10;	 rom[0][30][5] = 2'b11;	 rom[0][31][5] = 2'b11;	 rom[0][32][5] = 2'b10;	 rom[0][33][5] = 2'b00;	 rom[0][34][5] = 2'b00;	 rom[0][35][5] = 2'b00;	 rom[0][36][5] = 2'b00;	 rom[0][37][5] = 2'b00;	 rom[0][38][5] = 2'b00;	 rom[0][39][5] = 2'b00;
 rom[0][0][6] = 2'b00;	 rom[0][1][6] = 2'b00;	 rom[0][2][6] = 2'b00;	 rom[0][3][6] = 2'b00;	 rom[0][4][6] = 2'b00;	 rom[0][5][6] = 2'b00;	 rom[0][6][6] = 2'b00;	 rom[0][7][6] = 2'b00;	 rom[0][8][6] = 2'b00;	 rom[0][9][6] = 2'b00;	 rom[0][10][6] = 2'b00;	 rom[0][11][6] = 2'b00;	 rom[0][12][6] = 2'b00;	 rom[0][13][6] = 2'b00;	 rom[0][14][6] = 2'b00;	 rom[0][15][6] = 2'b00;	 rom[0][16][6] = 2'b00;	 rom[0][17][6] = 2'b00;	 rom[0][18][6] = 2'b00;	 rom[0][19][6] = 2'b10;	 rom[0][20][6] = 2'b10;	 rom[0][21][6] = 2'b10;	 rom[0][22][6] = 2'b10;	 rom[0][23][6] = 2'b10;	 rom[0][24][6] = 2'b10;	 rom[0][25][6] = 2'b00;	 rom[0][26][6] = 2'b00;	 rom[0][27][6] = 2'b00;	 rom[0][28][6] = 2'b00;	 rom[0][29][6] = 2'b10;	 rom[0][30][6] = 2'b11;	 rom[0][31][6] = 2'b11;	 rom[0][32][6] = 2'b10;	 rom[0][33][6] = 2'b00;	 rom[0][34][6] = 2'b00;	 rom[0][35][6] = 2'b00;	 rom[0][36][6] = 2'b00;	 rom[0][37][6] = 2'b00;	 rom[0][38][6] = 2'b00;	 rom[0][39][6] = 2'b00;
 rom[0][0][7] = 2'b00;	 rom[0][1][7] = 2'b00;	 rom[0][2][7] = 2'b00;	 rom[0][3][7] = 2'b00;	 rom[0][4][7] = 2'b00;	 rom[0][5][7] = 2'b00;	 rom[0][6][7] = 2'b00;	 rom[0][7][7] = 2'b00;	 rom[0][8][7] = 2'b00;	 rom[0][9][7] = 2'b10;	 rom[0][10][7] = 2'b10;	 rom[0][11][7] = 2'b10;	 rom[0][12][7] = 2'b10;	 rom[0][13][7] = 2'b10;	 rom[0][14][7] = 2'b10;	 rom[0][15][7] = 2'b00;	 rom[0][16][7] = 2'b00;	 rom[0][17][7] = 2'b00;	 rom[0][18][7] = 2'b10;	 rom[0][19][7] = 2'b10;	 rom[0][20][7] = 2'b11;	 rom[0][21][7] = 2'b11;	 rom[0][22][7] = 2'b11;	 rom[0][23][7] = 2'b11;	 rom[0][24][7] = 2'b10;	 rom[0][25][7] = 2'b10;	 rom[0][26][7] = 2'b00;	 rom[0][27][7] = 2'b00;	 rom[0][28][7] = 2'b00;	 rom[0][29][7] = 2'b10;	 rom[0][30][7] = 2'b11;	 rom[0][31][7] = 2'b11;	 rom[0][32][7] = 2'b10;	 rom[0][33][7] = 2'b00;	 rom[0][34][7] = 2'b00;	 rom[0][35][7] = 2'b00;	 rom[0][36][7] = 2'b00;	 rom[0][37][7] = 2'b00;	 rom[0][38][7] = 2'b00;	 rom[0][39][7] = 2'b00;
 rom[0][0][8] = 2'b00;	 rom[0][1][8] = 2'b00;	 rom[0][2][8] = 2'b00;	 rom[0][3][8] = 2'b00;	 rom[0][4][8] = 2'b00;	 rom[0][5][8] = 2'b00;	 rom[0][6][8] = 2'b00;	 rom[0][7][8] = 2'b00;	 rom[0][8][8] = 2'b10;	 rom[0][9][8] = 2'b10;	 rom[0][10][8] = 2'b11;	 rom[0][11][8] = 2'b11;	 rom[0][12][8] = 2'b11;	 rom[0][13][8] = 2'b11;	 rom[0][14][8] = 2'b10;	 rom[0][15][8] = 2'b10;	 rom[0][16][8] = 2'b00;	 rom[0][17][8] = 2'b00;	 rom[0][18][8] = 2'b10;	 rom[0][19][8] = 2'b11;	 rom[0][20][8] = 2'b11;	 rom[0][21][8] = 2'b11;	 rom[0][22][8] = 2'b11;	 rom[0][23][8] = 2'b11;	 rom[0][24][8] = 2'b11;	 rom[0][25][8] = 2'b10;	 rom[0][26][8] = 2'b10;	 rom[0][27][8] = 2'b00;	 rom[0][28][8] = 2'b00;	 rom[0][29][8] = 2'b10;	 rom[0][30][8] = 2'b11;	 rom[0][31][8] = 2'b11;	 rom[0][32][8] = 2'b10;	 rom[0][33][8] = 2'b10;	 rom[0][34][8] = 2'b00;	 rom[0][35][8] = 2'b00;	 rom[0][36][8] = 2'b00;	 rom[0][37][8] = 2'b00;	 rom[0][38][8] = 2'b00;	 rom[0][39][8] = 2'b00;
 rom[0][0][9] = 2'b00;	 rom[0][1][9] = 2'b00;	 rom[0][2][9] = 2'b00;	 rom[0][3][9] = 2'b00;	 rom[0][4][9] = 2'b00;	 rom[0][5][9] = 2'b00;	 rom[0][6][9] = 2'b00;	 rom[0][7][9] = 2'b10;	 rom[0][8][9] = 2'b10;	 rom[0][9][9] = 2'b11;	 rom[0][10][9] = 2'b11;	 rom[0][11][9] = 2'b11;	 rom[0][12][9] = 2'b11;	 rom[0][13][9] = 2'b11;	 rom[0][14][9] = 2'b11;	 rom[0][15][9] = 2'b10;	 rom[0][16][9] = 2'b10;	 rom[0][17][9] = 2'b00;	 rom[0][18][9] = 2'b10;	 rom[0][19][9] = 2'b11;	 rom[0][20][9] = 2'b11;	 rom[0][21][9] = 2'b11;	 rom[0][22][9] = 2'b11;	 rom[0][23][9] = 2'b11;	 rom[0][24][9] = 2'b11;	 rom[0][25][9] = 2'b11;	 rom[0][26][9] = 2'b10;	 rom[0][27][9] = 2'b00;	 rom[0][28][9] = 2'b00;	 rom[0][29][9] = 2'b10;	 rom[0][30][9] = 2'b11;	 rom[0][31][9] = 2'b11;	 rom[0][32][9] = 2'b10;	 rom[0][33][9] = 2'b10;	 rom[0][34][9] = 2'b10;	 rom[0][35][9] = 2'b00;	 rom[0][36][9] = 2'b00;	 rom[0][37][9] = 2'b00;	 rom[0][38][9] = 2'b00;	 rom[0][39][9] = 2'b00;
 rom[0][0][10] = 2'b00;	 rom[0][1][10] = 2'b00;	 rom[0][2][10] = 2'b00;	 rom[0][3][10] = 2'b00;	 rom[0][4][10] = 2'b00;	 rom[0][5][10] = 2'b00;	 rom[0][6][10] = 2'b00;	 rom[0][7][10] = 2'b10;	 rom[0][8][10] = 2'b11;	 rom[0][9][10] = 2'b11;	 rom[0][10][10] = 2'b11;	 rom[0][11][10] = 2'b11;	 rom[0][12][10] = 2'b11;	 rom[0][13][10] = 2'b11;	 rom[0][14][10] = 2'b10;	 rom[0][15][10] = 2'b10;	 rom[0][16][10] = 2'b10;	 rom[0][17][10] = 2'b10;	 rom[0][18][10] = 2'b10;	 rom[0][19][10] = 2'b10;	 rom[0][20][10] = 2'b10;	 rom[0][21][10] = 2'b10;	 rom[0][22][10] = 2'b10;	 rom[0][23][10] = 2'b10;	 rom[0][24][10] = 2'b10;	 rom[0][25][10] = 2'b10;	 rom[0][26][10] = 2'b10;	 rom[0][27][10] = 2'b00;	 rom[0][28][10] = 2'b00;	 rom[0][29][10] = 2'b10;	 rom[0][30][10] = 2'b11;	 rom[0][31][10] = 2'b11;	 rom[0][32][10] = 2'b10;	 rom[0][33][10] = 2'b01;	 rom[0][34][10] = 2'b10;	 rom[0][35][10] = 2'b00;	 rom[0][36][10] = 2'b00;	 rom[0][37][10] = 2'b00;	 rom[0][38][10] = 2'b00;	 rom[0][39][10] = 2'b00;
 rom[0][0][11] = 2'b00;	 rom[0][1][11] = 2'b00;	 rom[0][2][11] = 2'b00;	 rom[0][3][11] = 2'b00;	 rom[0][4][11] = 2'b00;	 rom[0][5][11] = 2'b00;	 rom[0][6][11] = 2'b00;	 rom[0][7][11] = 2'b10;	 rom[0][8][11] = 2'b11;	 rom[0][9][11] = 2'b11;	 rom[0][10][11] = 2'b11;	 rom[0][11][11] = 2'b11;	 rom[0][12][11] = 2'b10;	 rom[0][13][11] = 2'b10;	 rom[0][14][11] = 2'b10;	 rom[0][15][11] = 2'b10;	 rom[0][16][11] = 2'b10;	 rom[0][17][11] = 2'b10;	 rom[0][18][11] = 2'b10;	 rom[0][19][11] = 2'b10;	 rom[0][20][11] = 2'b10;	 rom[0][21][11] = 2'b10;	 rom[0][22][11] = 2'b10;	 rom[0][23][11] = 2'b10;	 rom[0][24][11] = 2'b10;	 rom[0][25][11] = 2'b10;	 rom[0][26][11] = 2'b10;	 rom[0][27][11] = 2'b10;	 rom[0][28][11] = 2'b00;	 rom[0][29][11] = 2'b10;	 rom[0][30][11] = 2'b11;	 rom[0][31][11] = 2'b11;	 rom[0][32][11] = 2'b10;	 rom[0][33][11] = 2'b01;	 rom[0][34][11] = 2'b10;	 rom[0][35][11] = 2'b10;	 rom[0][36][11] = 2'b10;	 rom[0][37][11] = 2'b10;	 rom[0][38][11] = 2'b10;	 rom[0][39][11] = 2'b10;
 rom[0][0][12] = 2'b00;	 rom[0][1][12] = 2'b00;	 rom[0][2][12] = 2'b00;	 rom[0][3][12] = 2'b00;	 rom[0][4][12] = 2'b00;	 rom[0][5][12] = 2'b00;	 rom[0][6][12] = 2'b00;	 rom[0][7][12] = 2'b10;	 rom[0][8][12] = 2'b11;	 rom[0][9][12] = 2'b11;	 rom[0][10][12] = 2'b11;	 rom[0][11][12] = 2'b11;	 rom[0][12][12] = 2'b10;	 rom[0][13][12] = 2'b10;	 rom[0][14][12] = 2'b01;	 rom[0][15][12] = 2'b01;	 rom[0][16][12] = 2'b01;	 rom[0][17][12] = 2'b01;	 rom[0][18][12] = 2'b01;	 rom[0][19][12] = 2'b01;	 rom[0][20][12] = 2'b01;	 rom[0][21][12] = 2'b01;	 rom[0][22][12] = 2'b01;	 rom[0][23][12] = 2'b01;	 rom[0][24][12] = 2'b01;	 rom[0][25][12] = 2'b01;	 rom[0][26][12] = 2'b10;	 rom[0][27][12] = 2'b10;	 rom[0][28][12] = 2'b00;	 rom[0][29][12] = 2'b10;	 rom[0][30][12] = 2'b11;	 rom[0][31][12] = 2'b11;	 rom[0][32][12] = 2'b10;	 rom[0][33][12] = 2'b01;	 rom[0][34][12] = 2'b01;	 rom[0][35][12] = 2'b10;	 rom[0][36][12] = 2'b10;	 rom[0][37][12] = 2'b11;	 rom[0][38][12] = 2'b11;	 rom[0][39][12] = 2'b10;
 rom[0][0][13] = 2'b00;	 rom[0][1][13] = 2'b00;	 rom[0][2][13] = 2'b00;	 rom[0][3][13] = 2'b00;	 rom[0][4][13] = 2'b00;	 rom[0][5][13] = 2'b00;	 rom[0][6][13] = 2'b00;	 rom[0][7][13] = 2'b10;	 rom[0][8][13] = 2'b11;	 rom[0][9][13] = 2'b11;	 rom[0][10][13] = 2'b10;	 rom[0][11][13] = 2'b10;	 rom[0][12][13] = 2'b10;	 rom[0][13][13] = 2'b01;	 rom[0][14][13] = 2'b01;	 rom[0][15][13] = 2'b01;	 rom[0][16][13] = 2'b01;	 rom[0][17][13] = 2'b01;	 rom[0][18][13] = 2'b01;	 rom[0][19][13] = 2'b01;	 rom[0][20][13] = 2'b01;	 rom[0][21][13] = 2'b01;	 rom[0][22][13] = 2'b01;	 rom[0][23][13] = 2'b01;	 rom[0][24][13] = 2'b01;	 rom[0][25][13] = 2'b01;	 rom[0][26][13] = 2'b01;	 rom[0][27][13] = 2'b10;	 rom[0][28][13] = 2'b10;	 rom[0][29][13] = 2'b10;	 rom[0][30][13] = 2'b11;	 rom[0][31][13] = 2'b11;	 rom[0][32][13] = 2'b10;	 rom[0][33][13] = 2'b01;	 rom[0][34][13] = 2'b01;	 rom[0][35][13] = 2'b01;	 rom[0][36][13] = 2'b10;	 rom[0][37][13] = 2'b11;	 rom[0][38][13] = 2'b11;	 rom[0][39][13] = 2'b10;
 rom[0][0][14] = 2'b00;	 rom[0][1][14] = 2'b00;	 rom[0][2][14] = 2'b00;	 rom[0][3][14] = 2'b00;	 rom[0][4][14] = 2'b00;	 rom[0][5][14] = 2'b00;	 rom[0][6][14] = 2'b00;	 rom[0][7][14] = 2'b10;	 rom[0][8][14] = 2'b11;	 rom[0][9][14] = 2'b10;	 rom[0][10][14] = 2'b10;	 rom[0][11][14] = 2'b10;	 rom[0][12][14] = 2'b01;	 rom[0][13][14] = 2'b01;	 rom[0][14][14] = 2'b01;	 rom[0][15][14] = 2'b01;	 rom[0][16][14] = 2'b01;	 rom[0][17][14] = 2'b01;	 rom[0][18][14] = 2'b01;	 rom[0][19][14] = 2'b01;	 rom[0][20][14] = 2'b01;	 rom[0][21][14] = 2'b01;	 rom[0][22][14] = 2'b01;	 rom[0][23][14] = 2'b01;	 rom[0][24][14] = 2'b01;	 rom[0][25][14] = 2'b01;	 rom[0][26][14] = 2'b01;	 rom[0][27][14] = 2'b01;	 rom[0][28][14] = 2'b10;	 rom[0][29][14] = 2'b10;	 rom[0][30][14] = 2'b11;	 rom[0][31][14] = 2'b11;	 rom[0][32][14] = 2'b10;	 rom[0][33][14] = 2'b10;	 rom[0][34][14] = 2'b01;	 rom[0][35][14] = 2'b01;	 rom[0][36][14] = 2'b10;	 rom[0][37][14] = 2'b10;	 rom[0][38][14] = 2'b11;	 rom[0][39][14] = 2'b10;
 rom[0][0][15] = 2'b00;	 rom[0][1][15] = 2'b00;	 rom[0][2][15] = 2'b00;	 rom[0][3][15] = 2'b00;	 rom[0][4][15] = 2'b00;	 rom[0][5][15] = 2'b00;	 rom[0][6][15] = 2'b00;	 rom[0][7][15] = 2'b10;	 rom[0][8][15] = 2'b10;	 rom[0][9][15] = 2'b10;	 rom[0][10][15] = 2'b10;	 rom[0][11][15] = 2'b01;	 rom[0][12][15] = 2'b01;	 rom[0][13][15] = 2'b01;	 rom[0][14][15] = 2'b01;	 rom[0][15][15] = 2'b01;	 rom[0][16][15] = 2'b01;	 rom[0][17][15] = 2'b01;	 rom[0][18][15] = 2'b01;	 rom[0][19][15] = 2'b01;	 rom[0][20][15] = 2'b01;	 rom[0][21][15] = 2'b01;	 rom[0][22][15] = 2'b01;	 rom[0][23][15] = 2'b01;	 rom[0][24][15] = 2'b01;	 rom[0][25][15] = 2'b01;	 rom[0][26][15] = 2'b01;	 rom[0][27][15] = 2'b01;	 rom[0][28][15] = 2'b01;	 rom[0][29][15] = 2'b10;	 rom[0][30][15] = 2'b10;	 rom[0][31][15] = 2'b11;	 rom[0][32][15] = 2'b10;	 rom[0][33][15] = 2'b10;	 rom[0][34][15] = 2'b01;	 rom[0][35][15] = 2'b01;	 rom[0][36][15] = 2'b01;	 rom[0][37][15] = 2'b10;	 rom[0][38][15] = 2'b10;	 rom[0][39][15] = 2'b10;
 rom[0][0][16] = 2'b00;	 rom[0][1][16] = 2'b00;	 rom[0][2][16] = 2'b00;	 rom[0][3][16] = 2'b00;	 rom[0][4][16] = 2'b00;	 rom[0][5][16] = 2'b00;	 rom[0][6][16] = 2'b00;	 rom[0][7][16] = 2'b00;	 rom[0][8][16] = 2'b10;	 rom[0][9][16] = 2'b10;	 rom[0][10][16] = 2'b01;	 rom[0][11][16] = 2'b01;	 rom[0][12][16] = 2'b01;	 rom[0][13][16] = 2'b01;	 rom[0][14][16] = 2'b01;	 rom[0][15][16] = 2'b01;	 rom[0][16][16] = 2'b01;	 rom[0][17][16] = 2'b01;	 rom[0][18][16] = 2'b01;	 rom[0][19][16] = 2'b01;	 rom[0][20][16] = 2'b01;	 rom[0][21][16] = 2'b01;	 rom[0][22][16] = 2'b01;	 rom[0][23][16] = 2'b01;	 rom[0][24][16] = 2'b01;	 rom[0][25][16] = 2'b01;	 rom[0][26][16] = 2'b01;	 rom[0][27][16] = 2'b01;	 rom[0][28][16] = 2'b01;	 rom[0][29][16] = 2'b01;	 rom[0][30][16] = 2'b10;	 rom[0][31][16] = 2'b10;	 rom[0][32][16] = 2'b10;	 rom[0][33][16] = 2'b10;	 rom[0][34][16] = 2'b01;	 rom[0][35][16] = 2'b01;	 rom[0][36][16] = 2'b01;	 rom[0][37][16] = 2'b10;	 rom[0][38][16] = 2'b00;	 rom[0][39][16] = 2'b00;
 rom[0][0][17] = 2'b00;	 rom[0][1][17] = 2'b00;	 rom[0][2][17] = 2'b00;	 rom[0][3][17] = 2'b00;	 rom[0][4][17] = 2'b00;	 rom[0][5][17] = 2'b00;	 rom[0][6][17] = 2'b10;	 rom[0][7][17] = 2'b10;	 rom[0][8][17] = 2'b10;	 rom[0][9][17] = 2'b01;	 rom[0][10][17] = 2'b01;	 rom[0][11][17] = 2'b01;	 rom[0][12][17] = 2'b01;	 rom[0][13][17] = 2'b01;	 rom[0][14][17] = 2'b01;	 rom[0][15][17] = 2'b01;	 rom[0][16][17] = 2'b01;	 rom[0][17][17] = 2'b01;	 rom[0][18][17] = 2'b01;	 rom[0][19][17] = 2'b01;	 rom[0][20][17] = 2'b01;	 rom[0][21][17] = 2'b01;	 rom[0][22][17] = 2'b01;	 rom[0][23][17] = 2'b01;	 rom[0][24][17] = 2'b01;	 rom[0][25][17] = 2'b01;	 rom[0][26][17] = 2'b01;	 rom[0][27][17] = 2'b01;	 rom[0][28][17] = 2'b01;	 rom[0][29][17] = 2'b01;	 rom[0][30][17] = 2'b01;	 rom[0][31][17] = 2'b10;	 rom[0][32][17] = 2'b10;	 rom[0][33][17] = 2'b10;	 rom[0][34][17] = 2'b01;	 rom[0][35][17] = 2'b01;	 rom[0][36][17] = 2'b01;	 rom[0][37][17] = 2'b10;	 rom[0][38][17] = 2'b00;	 rom[0][39][17] = 2'b00;
 rom[0][0][18] = 2'b00;	 rom[0][1][18] = 2'b00;	 rom[0][2][18] = 2'b00;	 rom[0][3][18] = 2'b00;	 rom[0][4][18] = 2'b10;	 rom[0][5][18] = 2'b10;	 rom[0][6][18] = 2'b10;	 rom[0][7][18] = 2'b10;	 rom[0][8][18] = 2'b10;	 rom[0][9][18] = 2'b01;	 rom[0][10][18] = 2'b01;	 rom[0][11][18] = 2'b01;	 rom[0][12][18] = 2'b01;	 rom[0][13][18] = 2'b01;	 rom[0][14][18] = 2'b01;	 rom[0][15][18] = 2'b01;	 rom[0][16][18] = 2'b01;	 rom[0][17][18] = 2'b01;	 rom[0][18][18] = 2'b01;	 rom[0][19][18] = 2'b01;	 rom[0][20][18] = 2'b01;	 rom[0][21][18] = 2'b01;	 rom[0][22][18] = 2'b01;	 rom[0][23][18] = 2'b01;	 rom[0][24][18] = 2'b01;	 rom[0][25][18] = 2'b01;	 rom[0][26][18] = 2'b01;	 rom[0][27][18] = 2'b01;	 rom[0][28][18] = 2'b01;	 rom[0][29][18] = 2'b01;	 rom[0][30][18] = 2'b01;	 rom[0][31][18] = 2'b10;	 rom[0][32][18] = 2'b10;	 rom[0][33][18] = 2'b10;	 rom[0][34][18] = 2'b01;	 rom[0][35][18] = 2'b01;	 rom[0][36][18] = 2'b01;	 rom[0][37][18] = 2'b10;	 rom[0][38][18] = 2'b00;	 rom[0][39][18] = 2'b00;
 rom[0][0][19] = 2'b00;	 rom[0][1][19] = 2'b00;	 rom[0][2][19] = 2'b10;	 rom[0][3][19] = 2'b10;	 rom[0][4][19] = 2'b10;	 rom[0][5][19] = 2'b01;	 rom[0][6][19] = 2'b10;	 rom[0][7][19] = 2'b10;	 rom[0][8][19] = 2'b10;	 rom[0][9][19] = 2'b01;	 rom[0][10][19] = 2'b01;	 rom[0][11][19] = 2'b01;	 rom[0][12][19] = 2'b01;	 rom[0][13][19] = 2'b01;	 rom[0][14][19] = 2'b01;	 rom[0][15][19] = 2'b01;	 rom[0][16][19] = 2'b01;	 rom[0][17][19] = 2'b01;	 rom[0][18][19] = 2'b01;	 rom[0][19][19] = 2'b01;	 rom[0][20][19] = 2'b01;	 rom[0][21][19] = 2'b01;	 rom[0][22][19] = 2'b01;	 rom[0][23][19] = 2'b01;	 rom[0][24][19] = 2'b01;	 rom[0][25][19] = 2'b01;	 rom[0][26][19] = 2'b01;	 rom[0][27][19] = 2'b01;	 rom[0][28][19] = 2'b01;	 rom[0][29][19] = 2'b01;	 rom[0][30][19] = 2'b01;	 rom[0][31][19] = 2'b10;	 rom[0][32][19] = 2'b10;	 rom[0][33][19] = 2'b10;	 rom[0][34][19] = 2'b01;	 rom[0][35][19] = 2'b01;	 rom[0][36][19] = 2'b01;	 rom[0][37][19] = 2'b10;	 rom[0][38][19] = 2'b00;	 rom[0][39][19] = 2'b00;
 rom[0][0][20] = 2'b00;	 rom[0][1][20] = 2'b00;	 rom[0][2][20] = 2'b10;	 rom[0][3][20] = 2'b10;	 rom[0][4][20] = 2'b01;	 rom[0][5][20] = 2'b01;	 rom[0][6][20] = 2'b10;	 rom[0][7][20] = 2'b10;	 rom[0][8][20] = 2'b01;	 rom[0][9][20] = 2'b01;	 rom[0][10][20] = 2'b01;	 rom[0][11][20] = 2'b01;	 rom[0][12][20] = 2'b01;	 rom[0][13][20] = 2'b01;	 rom[0][14][20] = 2'b01;	 rom[0][15][20] = 2'b01;	 rom[0][16][20] = 2'b01;	 rom[0][17][20] = 2'b01;	 rom[0][18][20] = 2'b01;	 rom[0][19][20] = 2'b01;	 rom[0][20][20] = 2'b01;	 rom[0][21][20] = 2'b01;	 rom[0][22][20] = 2'b01;	 rom[0][23][20] = 2'b01;	 rom[0][24][20] = 2'b01;	 rom[0][25][20] = 2'b01;	 rom[0][26][20] = 2'b01;	 rom[0][27][20] = 2'b01;	 rom[0][28][20] = 2'b01;	 rom[0][29][20] = 2'b01;	 rom[0][30][20] = 2'b01;	 rom[0][31][20] = 2'b01;	 rom[0][32][20] = 2'b10;	 rom[0][33][20] = 2'b10;	 rom[0][34][20] = 2'b01;	 rom[0][35][20] = 2'b01;	 rom[0][36][20] = 2'b01;	 rom[0][37][20] = 2'b10;	 rom[0][38][20] = 2'b00;	 rom[0][39][20] = 2'b00;
 rom[0][0][21] = 2'b00;	 rom[0][1][21] = 2'b00;	 rom[0][2][21] = 2'b10;	 rom[0][3][21] = 2'b01;	 rom[0][4][21] = 2'b01;	 rom[0][5][21] = 2'b01;	 rom[0][6][21] = 2'b10;	 rom[0][7][21] = 2'b10;	 rom[0][8][21] = 2'b01;	 rom[0][9][21] = 2'b01;	 rom[0][10][21] = 2'b01;	 rom[0][11][21] = 2'b01;	 rom[0][12][21] = 2'b01;	 rom[0][13][21] = 2'b01;	 rom[0][14][21] = 2'b01;	 rom[0][15][21] = 2'b01;	 rom[0][16][21] = 2'b01;	 rom[0][17][21] = 2'b01;	 rom[0][18][21] = 2'b01;	 rom[0][19][21] = 2'b01;	 rom[0][20][21] = 2'b01;	 rom[0][21][21] = 2'b01;	 rom[0][22][21] = 2'b01;	 rom[0][23][21] = 2'b01;	 rom[0][24][21] = 2'b01;	 rom[0][25][21] = 2'b01;	 rom[0][26][21] = 2'b01;	 rom[0][27][21] = 2'b01;	 rom[0][28][21] = 2'b01;	 rom[0][29][21] = 2'b01;	 rom[0][30][21] = 2'b01;	 rom[0][31][21] = 2'b01;	 rom[0][32][21] = 2'b10;	 rom[0][33][21] = 2'b10;	 rom[0][34][21] = 2'b01;	 rom[0][35][21] = 2'b01;	 rom[0][36][21] = 2'b01;	 rom[0][37][21] = 2'b10;	 rom[0][38][21] = 2'b00;	 rom[0][39][21] = 2'b00;
 rom[0][0][22] = 2'b00;	 rom[0][1][22] = 2'b00;	 rom[0][2][22] = 2'b10;	 rom[0][3][22] = 2'b01;	 rom[0][4][22] = 2'b01;	 rom[0][5][22] = 2'b01;	 rom[0][6][22] = 2'b10;	 rom[0][7][22] = 2'b10;	 rom[0][8][22] = 2'b01;	 rom[0][9][22] = 2'b01;	 rom[0][10][22] = 2'b01;	 rom[0][11][22] = 2'b01;	 rom[0][12][22] = 2'b01;	 rom[0][13][22] = 2'b01;	 rom[0][14][22] = 2'b01;	 rom[0][15][22] = 2'b01;	 rom[0][16][22] = 2'b01;	 rom[0][17][22] = 2'b01;	 rom[0][18][22] = 2'b01;	 rom[0][19][22] = 2'b01;	 rom[0][20][22] = 2'b01;	 rom[0][21][22] = 2'b01;	 rom[0][22][22] = 2'b01;	 rom[0][23][22] = 2'b01;	 rom[0][24][22] = 2'b01;	 rom[0][25][22] = 2'b01;	 rom[0][26][22] = 2'b01;	 rom[0][27][22] = 2'b01;	 rom[0][28][22] = 2'b01;	 rom[0][29][22] = 2'b01;	 rom[0][30][22] = 2'b01;	 rom[0][31][22] = 2'b10;	 rom[0][32][22] = 2'b10;	 rom[0][33][22] = 2'b10;	 rom[0][34][22] = 2'b01;	 rom[0][35][22] = 2'b01;	 rom[0][36][22] = 2'b01;	 rom[0][37][22] = 2'b10;	 rom[0][38][22] = 2'b00;	 rom[0][39][22] = 2'b00;
 rom[0][0][23] = 2'b00;	 rom[0][1][23] = 2'b00;	 rom[0][2][23] = 2'b10;	 rom[0][3][23] = 2'b01;	 rom[0][4][23] = 2'b01;	 rom[0][5][23] = 2'b01;	 rom[0][6][23] = 2'b10;	 rom[0][7][23] = 2'b10;	 rom[0][8][23] = 2'b01;	 rom[0][9][23] = 2'b01;	 rom[0][10][23] = 2'b01;	 rom[0][11][23] = 2'b01;	 rom[0][12][23] = 2'b01;	 rom[0][13][23] = 2'b01;	 rom[0][14][23] = 2'b01;	 rom[0][15][23] = 2'b01;	 rom[0][16][23] = 2'b01;	 rom[0][17][23] = 2'b01;	 rom[0][18][23] = 2'b01;	 rom[0][19][23] = 2'b01;	 rom[0][20][23] = 2'b01;	 rom[0][21][23] = 2'b01;	 rom[0][22][23] = 2'b01;	 rom[0][23][23] = 2'b01;	 rom[0][24][23] = 2'b01;	 rom[0][25][23] = 2'b01;	 rom[0][26][23] = 2'b01;	 rom[0][27][23] = 2'b01;	 rom[0][28][23] = 2'b01;	 rom[0][29][23] = 2'b01;	 rom[0][30][23] = 2'b01;	 rom[0][31][23] = 2'b01;	 rom[0][32][23] = 2'b10;	 rom[0][33][23] = 2'b10;	 rom[0][34][23] = 2'b01;	 rom[0][35][23] = 2'b01;	 rom[0][36][23] = 2'b01;	 rom[0][37][23] = 2'b10;	 rom[0][38][23] = 2'b00;	 rom[0][39][23] = 2'b00;
 rom[0][0][24] = 2'b00;	 rom[0][1][24] = 2'b00;	 rom[0][2][24] = 2'b10;	 rom[0][3][24] = 2'b01;	 rom[0][4][24] = 2'b01;	 rom[0][5][24] = 2'b01;	 rom[0][6][24] = 2'b10;	 rom[0][7][24] = 2'b10;	 rom[0][8][24] = 2'b01;	 rom[0][9][24] = 2'b01;	 rom[0][10][24] = 2'b01;	 rom[0][11][24] = 2'b01;	 rom[0][12][24] = 2'b01;	 rom[0][13][24] = 2'b01;	 rom[0][14][24] = 2'b01;	 rom[0][15][24] = 2'b01;	 rom[0][16][24] = 2'b01;	 rom[0][17][24] = 2'b01;	 rom[0][18][24] = 2'b01;	 rom[0][19][24] = 2'b01;	 rom[0][20][24] = 2'b01;	 rom[0][21][24] = 2'b01;	 rom[0][22][24] = 2'b01;	 rom[0][23][24] = 2'b01;	 rom[0][24][24] = 2'b01;	 rom[0][25][24] = 2'b01;	 rom[0][26][24] = 2'b01;	 rom[0][27][24] = 2'b01;	 rom[0][28][24] = 2'b01;	 rom[0][29][24] = 2'b01;	 rom[0][30][24] = 2'b01;	 rom[0][31][24] = 2'b01;	 rom[0][32][24] = 2'b10;	 rom[0][33][24] = 2'b10;	 rom[0][34][24] = 2'b01;	 rom[0][35][24] = 2'b01;	 rom[0][36][24] = 2'b01;	 rom[0][37][24] = 2'b10;	 rom[0][38][24] = 2'b00;	 rom[0][39][24] = 2'b00;
 rom[0][0][25] = 2'b00;	 rom[0][1][25] = 2'b00;	 rom[0][2][25] = 2'b10;	 rom[0][3][25] = 2'b01;	 rom[0][4][25] = 2'b01;	 rom[0][5][25] = 2'b01;	 rom[0][6][25] = 2'b10;	 rom[0][7][25] = 2'b10;	 rom[0][8][25] = 2'b01;	 rom[0][9][25] = 2'b01;	 rom[0][10][25] = 2'b01;	 rom[0][11][25] = 2'b01;	 rom[0][12][25] = 2'b01;	 rom[0][13][25] = 2'b01;	 rom[0][14][25] = 2'b01;	 rom[0][15][25] = 2'b01;	 rom[0][16][25] = 2'b01;	 rom[0][17][25] = 2'b01;	 rom[0][18][25] = 2'b01;	 rom[0][19][25] = 2'b01;	 rom[0][20][25] = 2'b01;	 rom[0][21][25] = 2'b01;	 rom[0][22][25] = 2'b01;	 rom[0][23][25] = 2'b01;	 rom[0][24][25] = 2'b01;	 rom[0][25][25] = 2'b01;	 rom[0][26][25] = 2'b01;	 rom[0][27][25] = 2'b01;	 rom[0][28][25] = 2'b01;	 rom[0][29][25] = 2'b01;	 rom[0][30][25] = 2'b01;	 rom[0][31][25] = 2'b10;	 rom[0][32][25] = 2'b10;	 rom[0][33][25] = 2'b10;	 rom[0][34][25] = 2'b01;	 rom[0][35][25] = 2'b01;	 rom[0][36][25] = 2'b01;	 rom[0][37][25] = 2'b10;	 rom[0][38][25] = 2'b00;	 rom[0][39][25] = 2'b00;
 rom[0][0][26] = 2'b00;	 rom[0][1][26] = 2'b00;	 rom[0][2][26] = 2'b10;	 rom[0][3][26] = 2'b01;	 rom[0][4][26] = 2'b01;	 rom[0][5][26] = 2'b01;	 rom[0][6][26] = 2'b10;	 rom[0][7][26] = 2'b10;	 rom[0][8][26] = 2'b10;	 rom[0][9][26] = 2'b01;	 rom[0][10][26] = 2'b01;	 rom[0][11][26] = 2'b01;	 rom[0][12][26] = 2'b01;	 rom[0][13][26] = 2'b01;	 rom[0][14][26] = 2'b01;	 rom[0][15][26] = 2'b01;	 rom[0][16][26] = 2'b01;	 rom[0][17][26] = 2'b01;	 rom[0][18][26] = 2'b01;	 rom[0][19][26] = 2'b01;	 rom[0][20][26] = 2'b01;	 rom[0][21][26] = 2'b01;	 rom[0][22][26] = 2'b01;	 rom[0][23][26] = 2'b01;	 rom[0][24][26] = 2'b01;	 rom[0][25][26] = 2'b01;	 rom[0][26][26] = 2'b01;	 rom[0][27][26] = 2'b01;	 rom[0][28][26] = 2'b01;	 rom[0][29][26] = 2'b01;	 rom[0][30][26] = 2'b01;	 rom[0][31][26] = 2'b10;	 rom[0][32][26] = 2'b10;	 rom[0][33][26] = 2'b10;	 rom[0][34][26] = 2'b01;	 rom[0][35][26] = 2'b01;	 rom[0][36][26] = 2'b01;	 rom[0][37][26] = 2'b10;	 rom[0][38][26] = 2'b00;	 rom[0][39][26] = 2'b00;
 rom[0][0][27] = 2'b00;	 rom[0][1][27] = 2'b00;	 rom[0][2][27] = 2'b10;	 rom[0][3][27] = 2'b01;	 rom[0][4][27] = 2'b01;	 rom[0][5][27] = 2'b01;	 rom[0][6][27] = 2'b01;	 rom[0][7][27] = 2'b10;	 rom[0][8][27] = 2'b10;	 rom[0][9][27] = 2'b10;	 rom[0][10][27] = 2'b01;	 rom[0][11][27] = 2'b01;	 rom[0][12][27] = 2'b01;	 rom[0][13][27] = 2'b01;	 rom[0][14][27] = 2'b01;	 rom[0][15][27] = 2'b01;	 rom[0][16][27] = 2'b01;	 rom[0][17][27] = 2'b01;	 rom[0][18][27] = 2'b01;	 rom[0][19][27] = 2'b01;	 rom[0][20][27] = 2'b01;	 rom[0][21][27] = 2'b01;	 rom[0][22][27] = 2'b01;	 rom[0][23][27] = 2'b01;	 rom[0][24][27] = 2'b01;	 rom[0][25][27] = 2'b01;	 rom[0][26][27] = 2'b01;	 rom[0][27][27] = 2'b01;	 rom[0][28][27] = 2'b01;	 rom[0][29][27] = 2'b01;	 rom[0][30][27] = 2'b10;	 rom[0][31][27] = 2'b10;	 rom[0][32][27] = 2'b10;	 rom[0][33][27] = 2'b01;	 rom[0][34][27] = 2'b01;	 rom[0][35][27] = 2'b01;	 rom[0][36][27] = 2'b01;	 rom[0][37][27] = 2'b10;	 rom[0][38][27] = 2'b00;	 rom[0][39][27] = 2'b00;
 rom[0][0][28] = 2'b00;	 rom[0][1][28] = 2'b00;	 rom[0][2][28] = 2'b10;	 rom[0][3][28] = 2'b10;	 rom[0][4][28] = 2'b01;	 rom[0][5][28] = 2'b01;	 rom[0][6][28] = 2'b01;	 rom[0][7][28] = 2'b01;	 rom[0][8][28] = 2'b10;	 rom[0][9][28] = 2'b10;	 rom[0][10][28] = 2'b10;	 rom[0][11][28] = 2'b01;	 rom[0][12][28] = 2'b01;	 rom[0][13][28] = 2'b01;	 rom[0][14][28] = 2'b01;	 rom[0][15][28] = 2'b01;	 rom[0][16][28] = 2'b01;	 rom[0][17][28] = 2'b01;	 rom[0][18][28] = 2'b01;	 rom[0][19][28] = 2'b01;	 rom[0][20][28] = 2'b01;	 rom[0][21][28] = 2'b01;	 rom[0][22][28] = 2'b01;	 rom[0][23][28] = 2'b01;	 rom[0][24][28] = 2'b01;	 rom[0][25][28] = 2'b01;	 rom[0][26][28] = 2'b01;	 rom[0][27][28] = 2'b01;	 rom[0][28][28] = 2'b01;	 rom[0][29][28] = 2'b10;	 rom[0][30][28] = 2'b10;	 rom[0][31][28] = 2'b10;	 rom[0][32][28] = 2'b01;	 rom[0][33][28] = 2'b01;	 rom[0][34][28] = 2'b01;	 rom[0][35][28] = 2'b01;	 rom[0][36][28] = 2'b10;	 rom[0][37][28] = 2'b10;	 rom[0][38][28] = 2'b00;	 rom[0][39][28] = 2'b00;
 rom[0][0][29] = 2'b00;	 rom[0][1][29] = 2'b00;	 rom[0][2][29] = 2'b00;	 rom[0][3][29] = 2'b10;	 rom[0][4][29] = 2'b10;	 rom[0][5][29] = 2'b10;	 rom[0][6][29] = 2'b10;	 rom[0][7][29] = 2'b10;	 rom[0][8][29] = 2'b10;	 rom[0][9][29] = 2'b10;	 rom[0][10][29] = 2'b10;	 rom[0][11][29] = 2'b10;	 rom[0][12][29] = 2'b01;	 rom[0][13][29] = 2'b01;	 rom[0][14][29] = 2'b01;	 rom[0][15][29] = 2'b01;	 rom[0][16][29] = 2'b01;	 rom[0][17][29] = 2'b01;	 rom[0][18][29] = 2'b01;	 rom[0][19][29] = 2'b01;	 rom[0][20][29] = 2'b01;	 rom[0][21][29] = 2'b01;	 rom[0][22][29] = 2'b01;	 rom[0][23][29] = 2'b01;	 rom[0][24][29] = 2'b01;	 rom[0][25][29] = 2'b01;	 rom[0][26][29] = 2'b01;	 rom[0][27][29] = 2'b01;	 rom[0][28][29] = 2'b10;	 rom[0][29][29] = 2'b10;	 rom[0][30][29] = 2'b10;	 rom[0][31][29] = 2'b10;	 rom[0][32][29] = 2'b10;	 rom[0][33][29] = 2'b10;	 rom[0][34][29] = 2'b10;	 rom[0][35][29] = 2'b10;	 rom[0][36][29] = 2'b10;	 rom[0][37][29] = 2'b00;	 rom[0][38][29] = 2'b00;	 rom[0][39][29] = 2'b00;
 rom[0][0][30] = 2'b00;	 rom[0][1][30] = 2'b00;	 rom[0][2][30] = 2'b00;	 rom[0][3][30] = 2'b00;	 rom[0][4][30] = 2'b10;	 rom[0][5][30] = 2'b10;	 rom[0][6][30] = 2'b10;	 rom[0][7][30] = 2'b10;	 rom[0][8][30] = 2'b10;	 rom[0][9][30] = 2'b10;	 rom[0][10][30] = 2'b10;	 rom[0][11][30] = 2'b10;	 rom[0][12][30] = 2'b10;	 rom[0][13][30] = 2'b10;	 rom[0][14][30] = 2'b10;	 rom[0][15][30] = 2'b10;	 rom[0][16][30] = 2'b01;	 rom[0][17][30] = 2'b01;	 rom[0][18][30] = 2'b01;	 rom[0][19][30] = 2'b01;	 rom[0][20][30] = 2'b01;	 rom[0][21][30] = 2'b01;	 rom[0][22][30] = 2'b01;	 rom[0][23][30] = 2'b01;	 rom[0][24][30] = 2'b10;	 rom[0][25][30] = 2'b10;	 rom[0][26][30] = 2'b10;	 rom[0][27][30] = 2'b10;	 rom[0][28][30] = 2'b10;	 rom[0][29][30] = 2'b10;	 rom[0][30][30] = 2'b10;	 rom[0][31][30] = 2'b10;	 rom[0][32][30] = 2'b10;	 rom[0][33][30] = 2'b10;	 rom[0][34][30] = 2'b10;	 rom[0][35][30] = 2'b10;	 rom[0][36][30] = 2'b00;	 rom[0][37][30] = 2'b00;	 rom[0][38][30] = 2'b00;	 rom[0][39][30] = 2'b00;
 rom[0][0][31] = 2'b00;	 rom[0][1][31] = 2'b00;	 rom[0][2][31] = 2'b00;	 rom[0][3][31] = 2'b00;	 rom[0][4][31] = 2'b00;	 rom[0][5][31] = 2'b00;	 rom[0][6][31] = 2'b00;	 rom[0][7][31] = 2'b00;	 rom[0][8][31] = 2'b10;	 rom[0][9][31] = 2'b10;	 rom[0][10][31] = 2'b10;	 rom[0][11][31] = 2'b10;	 rom[0][12][31] = 2'b10;	 rom[0][13][31] = 2'b11;	 rom[0][14][31] = 2'b11;	 rom[0][15][31] = 2'b10;	 rom[0][16][31] = 2'b10;	 rom[0][17][31] = 2'b10;	 rom[0][18][31] = 2'b10;	 rom[0][19][31] = 2'b10;	 rom[0][20][31] = 2'b10;	 rom[0][21][31] = 2'b10;	 rom[0][22][31] = 2'b10;	 rom[0][23][31] = 2'b10;	 rom[0][24][31] = 2'b10;	 rom[0][25][31] = 2'b11;	 rom[0][26][31] = 2'b11;	 rom[0][27][31] = 2'b10;	 rom[0][28][31] = 2'b10;	 rom[0][29][31] = 2'b10;	 rom[0][30][31] = 2'b10;	 rom[0][31][31] = 2'b10;	 rom[0][32][31] = 2'b00;	 rom[0][33][31] = 2'b00;	 rom[0][34][31] = 2'b00;	 rom[0][35][31] = 2'b00;	 rom[0][36][31] = 2'b00;	 rom[0][37][31] = 2'b00;	 rom[0][38][31] = 2'b00;	 rom[0][39][31] = 2'b00;
 rom[0][0][32] = 2'b00;	 rom[0][1][32] = 2'b00;	 rom[0][2][32] = 2'b00;	 rom[0][3][32] = 2'b00;	 rom[0][4][32] = 2'b00;	 rom[0][5][32] = 2'b00;	 rom[0][6][32] = 2'b00;	 rom[0][7][32] = 2'b00;	 rom[0][8][32] = 2'b10;	 rom[0][9][32] = 2'b10;	 rom[0][10][32] = 2'b10;	 rom[0][11][32] = 2'b10;	 rom[0][12][32] = 2'b10;	 rom[0][13][32] = 2'b11;	 rom[0][14][32] = 2'b11;	 rom[0][15][32] = 2'b10;	 rom[0][16][32] = 2'b10;	 rom[0][17][32] = 2'b10;	 rom[0][18][32] = 2'b10;	 rom[0][19][32] = 2'b10;	 rom[0][20][32] = 2'b10;	 rom[0][21][32] = 2'b10;	 rom[0][22][32] = 2'b10;	 rom[0][23][32] = 2'b10;	 rom[0][24][32] = 2'b10;	 rom[0][25][32] = 2'b11;	 rom[0][26][32] = 2'b11;	 rom[0][27][32] = 2'b10;	 rom[0][28][32] = 2'b10;	 rom[0][29][32] = 2'b10;	 rom[0][30][32] = 2'b10;	 rom[0][31][32] = 2'b10;	 rom[0][32][32] = 2'b00;	 rom[0][33][32] = 2'b00;	 rom[0][34][32] = 2'b00;	 rom[0][35][32] = 2'b00;	 rom[0][36][32] = 2'b00;	 rom[0][37][32] = 2'b00;	 rom[0][38][32] = 2'b00;	 rom[0][39][32] = 2'b00;
 rom[0][0][33] = 2'b00;	 rom[0][1][33] = 2'b00;	 rom[0][2][33] = 2'b00;	 rom[0][3][33] = 2'b00;	 rom[0][4][33] = 2'b00;	 rom[0][5][33] = 2'b00;	 rom[0][6][33] = 2'b00;	 rom[0][7][33] = 2'b00;	 rom[0][8][33] = 2'b10;	 rom[0][9][33] = 2'b10;	 rom[0][10][33] = 2'b10;	 rom[0][11][33] = 2'b10;	 rom[0][12][33] = 2'b11;	 rom[0][13][33] = 2'b11;	 rom[0][14][33] = 2'b11;	 rom[0][15][33] = 2'b10;	 rom[0][16][33] = 2'b10;	 rom[0][17][33] = 2'b10;	 rom[0][18][33] = 2'b10;	 rom[0][19][33] = 2'b10;	 rom[0][20][33] = 2'b10;	 rom[0][21][33] = 2'b10;	 rom[0][22][33] = 2'b10;	 rom[0][23][33] = 2'b10;	 rom[0][24][33] = 2'b10;	 rom[0][25][33] = 2'b11;	 rom[0][26][33] = 2'b11;	 rom[0][27][33] = 2'b11;	 rom[0][28][33] = 2'b10;	 rom[0][29][33] = 2'b10;	 rom[0][30][33] = 2'b10;	 rom[0][31][33] = 2'b10;	 rom[0][32][33] = 2'b00;	 rom[0][33][33] = 2'b00;	 rom[0][34][33] = 2'b00;	 rom[0][35][33] = 2'b00;	 rom[0][36][33] = 2'b00;	 rom[0][37][33] = 2'b00;	 rom[0][38][33] = 2'b00;	 rom[0][39][33] = 2'b00;
 rom[0][0][34] = 2'b00;	 rom[0][1][34] = 2'b00;	 rom[0][2][34] = 2'b00;	 rom[0][3][34] = 2'b00;	 rom[0][4][34] = 2'b00;	 rom[0][5][34] = 2'b00;	 rom[0][6][34] = 2'b00;	 rom[0][7][34] = 2'b00;	 rom[0][8][34] = 2'b00;	 rom[0][9][34] = 2'b10;	 rom[0][10][34] = 2'b10;	 rom[0][11][34] = 2'b11;	 rom[0][12][34] = 2'b11;	 rom[0][13][34] = 2'b11;	 rom[0][14][34] = 2'b11;	 rom[0][15][34] = 2'b11;	 rom[0][16][34] = 2'b11;	 rom[0][17][34] = 2'b11;	 rom[0][18][34] = 2'b11;	 rom[0][19][34] = 2'b11;	 rom[0][20][34] = 2'b11;	 rom[0][21][34] = 2'b11;	 rom[0][22][34] = 2'b11;	 rom[0][23][34] = 2'b11;	 rom[0][24][34] = 2'b11;	 rom[0][25][34] = 2'b11;	 rom[0][26][34] = 2'b11;	 rom[0][27][34] = 2'b11;	 rom[0][28][34] = 2'b11;	 rom[0][29][34] = 2'b10;	 rom[0][30][34] = 2'b10;	 rom[0][31][34] = 2'b00;	 rom[0][32][34] = 2'b00;	 rom[0][33][34] = 2'b00;	 rom[0][34][34] = 2'b00;	 rom[0][35][34] = 2'b00;	 rom[0][36][34] = 2'b00;	 rom[0][37][34] = 2'b00;	 rom[0][38][34] = 2'b00;	 rom[0][39][34] = 2'b00;
 rom[0][0][35] = 2'b00;	 rom[0][1][35] = 2'b00;	 rom[0][2][35] = 2'b00;	 rom[0][3][35] = 2'b00;	 rom[0][4][35] = 2'b00;	 rom[0][5][35] = 2'b00;	 rom[0][6][35] = 2'b00;	 rom[0][7][35] = 2'b00;	 rom[0][8][35] = 2'b00;	 rom[0][9][35] = 2'b10;	 rom[0][10][35] = 2'b10;	 rom[0][11][35] = 2'b11;	 rom[0][12][35] = 2'b11;	 rom[0][13][35] = 2'b11;	 rom[0][14][35] = 2'b11;	 rom[0][15][35] = 2'b11;	 rom[0][16][35] = 2'b11;	 rom[0][17][35] = 2'b10;	 rom[0][18][35] = 2'b10;	 rom[0][19][35] = 2'b10;	 rom[0][20][35] = 2'b10;	 rom[0][21][35] = 2'b10;	 rom[0][22][35] = 2'b10;	 rom[0][23][35] = 2'b11;	 rom[0][24][35] = 2'b11;	 rom[0][25][35] = 2'b11;	 rom[0][26][35] = 2'b11;	 rom[0][27][35] = 2'b11;	 rom[0][28][35] = 2'b11;	 rom[0][29][35] = 2'b10;	 rom[0][30][35] = 2'b10;	 rom[0][31][35] = 2'b00;	 rom[0][32][35] = 2'b00;	 rom[0][33][35] = 2'b00;	 rom[0][34][35] = 2'b00;	 rom[0][35][35] = 2'b00;	 rom[0][36][35] = 2'b00;	 rom[0][37][35] = 2'b00;	 rom[0][38][35] = 2'b00;	 rom[0][39][35] = 2'b00;
 rom[0][0][36] = 2'b00;	 rom[0][1][36] = 2'b00;	 rom[0][2][36] = 2'b00;	 rom[0][3][36] = 2'b00;	 rom[0][4][36] = 2'b00;	 rom[0][5][36] = 2'b00;	 rom[0][6][36] = 2'b00;	 rom[0][7][36] = 2'b00;	 rom[0][8][36] = 2'b00;	 rom[0][9][36] = 2'b00;	 rom[0][10][36] = 2'b10;	 rom[0][11][36] = 2'b11;	 rom[0][12][36] = 2'b11;	 rom[0][13][36] = 2'b11;	 rom[0][14][36] = 2'b11;	 rom[0][15][36] = 2'b11;	 rom[0][16][36] = 2'b11;	 rom[0][17][36] = 2'b11;	 rom[0][18][36] = 2'b11;	 rom[0][19][36] = 2'b11;	 rom[0][20][36] = 2'b11;	 rom[0][21][36] = 2'b11;	 rom[0][22][36] = 2'b11;	 rom[0][23][36] = 2'b11;	 rom[0][24][36] = 2'b11;	 rom[0][25][36] = 2'b11;	 rom[0][26][36] = 2'b11;	 rom[0][27][36] = 2'b11;	 rom[0][28][36] = 2'b11;	 rom[0][29][36] = 2'b10;	 rom[0][30][36] = 2'b00;	 rom[0][31][36] = 2'b00;	 rom[0][32][36] = 2'b00;	 rom[0][33][36] = 2'b00;	 rom[0][34][36] = 2'b00;	 rom[0][35][36] = 2'b00;	 rom[0][36][36] = 2'b00;	 rom[0][37][36] = 2'b00;	 rom[0][38][36] = 2'b00;	 rom[0][39][36] = 2'b00;
 rom[0][0][37] = 2'b00;	 rom[0][1][37] = 2'b00;	 rom[0][2][37] = 2'b00;	 rom[0][3][37] = 2'b00;	 rom[0][4][37] = 2'b00;	 rom[0][5][37] = 2'b00;	 rom[0][6][37] = 2'b00;	 rom[0][7][37] = 2'b00;	 rom[0][8][37] = 2'b00;	 rom[0][9][37] = 2'b00;	 rom[0][10][37] = 2'b10;	 rom[0][11][37] = 2'b10;	 rom[0][12][37] = 2'b10;	 rom[0][13][37] = 2'b10;	 rom[0][14][37] = 2'b10;	 rom[0][15][37] = 2'b10;	 rom[0][16][37] = 2'b10;	 rom[0][17][37] = 2'b10;	 rom[0][18][37] = 2'b10;	 rom[0][19][37] = 2'b10;	 rom[0][20][37] = 2'b10;	 rom[0][21][37] = 2'b10;	 rom[0][22][37] = 2'b10;	 rom[0][23][37] = 2'b10;	 rom[0][24][37] = 2'b10;	 rom[0][25][37] = 2'b10;	 rom[0][26][37] = 2'b10;	 rom[0][27][37] = 2'b10;	 rom[0][28][37] = 2'b10;	 rom[0][29][37] = 2'b10;	 rom[0][30][37] = 2'b00;	 rom[0][31][37] = 2'b00;	 rom[0][32][37] = 2'b00;	 rom[0][33][37] = 2'b00;	 rom[0][34][37] = 2'b00;	 rom[0][35][37] = 2'b00;	 rom[0][36][37] = 2'b00;	 rom[0][37][37] = 2'b00;	 rom[0][38][37] = 2'b00;	 rom[0][39][37] = 2'b00;
 rom[0][0][38] = 2'b00;	 rom[0][1][38] = 2'b00;	 rom[0][2][38] = 2'b00;	 rom[0][3][38] = 2'b00;	 rom[0][4][38] = 2'b00;	 rom[0][5][38] = 2'b00;	 rom[0][6][38] = 2'b00;	 rom[0][7][38] = 2'b00;	 rom[0][8][38] = 2'b00;	 rom[0][9][38] = 2'b00;	 rom[0][10][38] = 2'b00;	 rom[0][11][38] = 2'b00;	 rom[0][12][38] = 2'b00;	 rom[0][13][38] = 2'b00;	 rom[0][14][38] = 2'b00;	 rom[0][15][38] = 2'b00;	 rom[0][16][38] = 2'b00;	 rom[0][17][38] = 2'b00;	 rom[0][18][38] = 2'b00;	 rom[0][19][38] = 2'b00;	 rom[0][20][38] = 2'b00;	 rom[0][21][38] = 2'b00;	 rom[0][22][38] = 2'b00;	 rom[0][23][38] = 2'b00;	 rom[0][24][38] = 2'b00;	 rom[0][25][38] = 2'b00;	 rom[0][26][38] = 2'b00;	 rom[0][27][38] = 2'b00;	 rom[0][28][38] = 2'b00;	 rom[0][29][38] = 2'b00;	 rom[0][30][38] = 2'b00;	 rom[0][31][38] = 2'b00;	 rom[0][32][38] = 2'b00;	 rom[0][33][38] = 2'b00;	 rom[0][34][38] = 2'b00;	 rom[0][35][38] = 2'b00;	 rom[0][36][38] = 2'b00;	 rom[0][37][38] = 2'b00;	 rom[0][38][38] = 2'b00;	 rom[0][39][38] = 2'b00;
 rom[0][0][39] = 2'b00;	 rom[0][1][39] = 2'b00;	 rom[0][2][39] = 2'b00;	 rom[0][3][39] = 2'b00;	 rom[0][4][39] = 2'b00;	 rom[0][5][39] = 2'b00;	 rom[0][6][39] = 2'b00;	 rom[0][7][39] = 2'b00;	 rom[0][8][39] = 2'b00;	 rom[0][9][39] = 2'b00;	 rom[0][10][39] = 2'b00;	 rom[0][11][39] = 2'b00;	 rom[0][12][39] = 2'b00;	 rom[0][13][39] = 2'b00;	 rom[0][14][39] = 2'b00;	 rom[0][15][39] = 2'b00;	 rom[0][16][39] = 2'b00;	 rom[0][17][39] = 2'b00;	 rom[0][18][39] = 2'b00;	 rom[0][19][39] = 2'b00;	 rom[0][20][39] = 2'b00;	 rom[0][21][39] = 2'b00;	 rom[0][22][39] = 2'b00;	 rom[0][23][39] = 2'b00;	 rom[0][24][39] = 2'b00;	 rom[0][25][39] = 2'b00;	 rom[0][26][39] = 2'b00;	 rom[0][27][39] = 2'b00;	 rom[0][28][39] = 2'b00;	 rom[0][29][39] = 2'b00;	 rom[0][30][39] = 2'b00;	 rom[0][31][39] = 2'b00;	 rom[0][32][39] = 2'b00;	 rom[0][33][39] = 2'b00;	 rom[0][34][39] = 2'b00;	 rom[0][35][39] = 2'b00;	 rom[0][36][39] = 2'b00;	 rom[0][37][39] = 2'b00;	 rom[0][38][39] = 2'b00;	 rom[0][39][39] = 2'b00;

 rom[1][0][0] = 2'b00;	 rom[1][1][0] = 2'b00;	 rom[1][2][0] = 2'b00;	 rom[1][3][0] = 2'b00;	 rom[1][4][0] = 2'b00;	 rom[1][5][0] = 2'b00;	 rom[1][6][0] = 2'b00;	 rom[1][7][0] = 2'b00;	 rom[1][8][0] = 2'b00;	 rom[1][9][0] = 2'b00;	 rom[1][10][0] = 2'b00;	 rom[1][11][0] = 2'b00;	 rom[1][12][0] = 2'b00;	 rom[1][13][0] = 2'b00;	 rom[1][14][0] = 2'b00;	 rom[1][15][0] = 2'b00;	 rom[1][16][0] = 2'b00;	 rom[1][17][0] = 2'b00;	 rom[1][18][0] = 2'b00;	 rom[1][19][0] = 2'b00;	 rom[1][20][0] = 2'b00;	 rom[1][21][0] = 2'b00;	 rom[1][22][0] = 2'b00;	 rom[1][23][0] = 2'b00;	 rom[1][24][0] = 2'b00;	 rom[1][25][0] = 2'b00;	 rom[1][26][0] = 2'b00;	 rom[1][27][0] = 2'b00;	 rom[1][28][0] = 2'b00;	 rom[1][29][0] = 2'b00;	 rom[1][30][0] = 2'b00;	 rom[1][31][0] = 2'b00;	 rom[1][32][0] = 2'b00;	 rom[1][33][0] = 2'b00;	 rom[1][34][0] = 2'b00;	 rom[1][35][0] = 2'b00;	 rom[1][36][0] = 2'b00;	 rom[1][37][0] = 2'b00;	 rom[1][38][0] = 2'b00;	 rom[1][39][0] = 2'b00;
 rom[1][0][1] = 2'b00;	 rom[1][1][1] = 2'b00;	 rom[1][2][1] = 2'b00;	 rom[1][3][1] = 2'b00;	 rom[1][4][1] = 2'b00;	 rom[1][5][1] = 2'b00;	 rom[1][6][1] = 2'b00;	 rom[1][7][1] = 2'b00;	 rom[1][8][1] = 2'b00;	 rom[1][9][1] = 2'b00;	 rom[1][10][1] = 2'b00;	 rom[1][11][1] = 2'b00;	 rom[1][12][1] = 2'b00;	 rom[1][13][1] = 2'b00;	 rom[1][14][1] = 2'b00;	 rom[1][15][1] = 2'b00;	 rom[1][16][1] = 2'b00;	 rom[1][17][1] = 2'b00;	 rom[1][18][1] = 2'b00;	 rom[1][19][1] = 2'b00;	 rom[1][20][1] = 2'b00;	 rom[1][21][1] = 2'b00;	 rom[1][22][1] = 2'b00;	 rom[1][23][1] = 2'b00;	 rom[1][24][1] = 2'b00;	 rom[1][25][1] = 2'b00;	 rom[1][26][1] = 2'b00;	 rom[1][27][1] = 2'b00;	 rom[1][28][1] = 2'b00;	 rom[1][29][1] = 2'b00;	 rom[1][30][1] = 2'b00;	 rom[1][31][1] = 2'b00;	 rom[1][32][1] = 2'b00;	 rom[1][33][1] = 2'b00;	 rom[1][34][1] = 2'b00;	 rom[1][35][1] = 2'b00;	 rom[1][36][1] = 2'b00;	 rom[1][37][1] = 2'b00;	 rom[1][38][1] = 2'b00;	 rom[1][39][1] = 2'b00;
 rom[1][0][2] = 2'b00;	 rom[1][1][2] = 2'b00;	 rom[1][2][2] = 2'b00;	 rom[1][3][2] = 2'b00;	 rom[1][4][2] = 2'b00;	 rom[1][5][2] = 2'b00;	 rom[1][6][2] = 2'b00;	 rom[1][7][2] = 2'b00;	 rom[1][8][2] = 2'b00;	 rom[1][9][2] = 2'b00;	 rom[1][10][2] = 2'b10;	 rom[1][11][2] = 2'b10;	 rom[1][12][2] = 2'b10;	 rom[1][13][2] = 2'b10;	 rom[1][14][2] = 2'b10;	 rom[1][15][2] = 2'b10;	 rom[1][16][2] = 2'b10;	 rom[1][17][2] = 2'b10;	 rom[1][18][2] = 2'b10;	 rom[1][19][2] = 2'b10;	 rom[1][20][2] = 2'b10;	 rom[1][21][2] = 2'b10;	 rom[1][22][2] = 2'b10;	 rom[1][23][2] = 2'b10;	 rom[1][24][2] = 2'b10;	 rom[1][25][2] = 2'b10;	 rom[1][26][2] = 2'b10;	 rom[1][27][2] = 2'b10;	 rom[1][28][2] = 2'b10;	 rom[1][29][2] = 2'b10;	 rom[1][30][2] = 2'b00;	 rom[1][31][2] = 2'b00;	 rom[1][32][2] = 2'b00;	 rom[1][33][2] = 2'b00;	 rom[1][34][2] = 2'b00;	 rom[1][35][2] = 2'b00;	 rom[1][36][2] = 2'b00;	 rom[1][37][2] = 2'b00;	 rom[1][38][2] = 2'b00;	 rom[1][39][2] = 2'b00;
 rom[1][0][3] = 2'b00;	 rom[1][1][3] = 2'b00;	 rom[1][2][3] = 2'b00;	 rom[1][3][3] = 2'b00;	 rom[1][4][3] = 2'b00;	 rom[1][5][3] = 2'b00;	 rom[1][6][3] = 2'b00;	 rom[1][7][3] = 2'b00;	 rom[1][8][3] = 2'b00;	 rom[1][9][3] = 2'b00;	 rom[1][10][3] = 2'b10;	 rom[1][11][3] = 2'b11;	 rom[1][12][3] = 2'b11;	 rom[1][13][3] = 2'b11;	 rom[1][14][3] = 2'b11;	 rom[1][15][3] = 2'b11;	 rom[1][16][3] = 2'b11;	 rom[1][17][3] = 2'b11;	 rom[1][18][3] = 2'b11;	 rom[1][19][3] = 2'b11;	 rom[1][20][3] = 2'b11;	 rom[1][21][3] = 2'b11;	 rom[1][22][3] = 2'b11;	 rom[1][23][3] = 2'b11;	 rom[1][24][3] = 2'b11;	 rom[1][25][3] = 2'b11;	 rom[1][26][3] = 2'b11;	 rom[1][27][3] = 2'b11;	 rom[1][28][3] = 2'b11;	 rom[1][29][3] = 2'b10;	 rom[1][30][3] = 2'b00;	 rom[1][31][3] = 2'b00;	 rom[1][32][3] = 2'b00;	 rom[1][33][3] = 2'b00;	 rom[1][34][3] = 2'b00;	 rom[1][35][3] = 2'b00;	 rom[1][36][3] = 2'b00;	 rom[1][37][3] = 2'b00;	 rom[1][38][3] = 2'b00;	 rom[1][39][3] = 2'b00;
 rom[1][0][4] = 2'b00;	 rom[1][1][4] = 2'b00;	 rom[1][2][4] = 2'b00;	 rom[1][3][4] = 2'b00;	 rom[1][4][4] = 2'b00;	 rom[1][5][4] = 2'b00;	 rom[1][6][4] = 2'b00;	 rom[1][7][4] = 2'b00;	 rom[1][8][4] = 2'b00;	 rom[1][9][4] = 2'b10;	 rom[1][10][4] = 2'b10;	 rom[1][11][4] = 2'b11;	 rom[1][12][4] = 2'b11;	 rom[1][13][4] = 2'b11;	 rom[1][14][4] = 2'b11;	 rom[1][15][4] = 2'b11;	 rom[1][16][4] = 2'b11;	 rom[1][17][4] = 2'b10;	 rom[1][18][4] = 2'b10;	 rom[1][19][4] = 2'b10;	 rom[1][20][4] = 2'b10;	 rom[1][21][4] = 2'b10;	 rom[1][22][4] = 2'b10;	 rom[1][23][4] = 2'b11;	 rom[1][24][4] = 2'b11;	 rom[1][25][4] = 2'b11;	 rom[1][26][4] = 2'b11;	 rom[1][27][4] = 2'b11;	 rom[1][28][4] = 2'b11;	 rom[1][29][4] = 2'b10;	 rom[1][30][4] = 2'b10;	 rom[1][31][4] = 2'b00;	 rom[1][32][4] = 2'b00;	 rom[1][33][4] = 2'b00;	 rom[1][34][4] = 2'b00;	 rom[1][35][4] = 2'b00;	 rom[1][36][4] = 2'b00;	 rom[1][37][4] = 2'b00;	 rom[1][38][4] = 2'b00;	 rom[1][39][4] = 2'b00;
 rom[1][0][5] = 2'b00;	 rom[1][1][5] = 2'b00;	 rom[1][2][5] = 2'b00;	 rom[1][3][5] = 2'b00;	 rom[1][4][5] = 2'b00;	 rom[1][5][5] = 2'b00;	 rom[1][6][5] = 2'b00;	 rom[1][7][5] = 2'b00;	 rom[1][8][5] = 2'b00;	 rom[1][9][5] = 2'b10;	 rom[1][10][5] = 2'b10;	 rom[1][11][5] = 2'b11;	 rom[1][12][5] = 2'b11;	 rom[1][13][5] = 2'b11;	 rom[1][14][5] = 2'b11;	 rom[1][15][5] = 2'b11;	 rom[1][16][5] = 2'b11;	 rom[1][17][5] = 2'b11;	 rom[1][18][5] = 2'b11;	 rom[1][19][5] = 2'b11;	 rom[1][20][5] = 2'b11;	 rom[1][21][5] = 2'b11;	 rom[1][22][5] = 2'b11;	 rom[1][23][5] = 2'b11;	 rom[1][24][5] = 2'b11;	 rom[1][25][5] = 2'b11;	 rom[1][26][5] = 2'b11;	 rom[1][27][5] = 2'b11;	 rom[1][28][5] = 2'b11;	 rom[1][29][5] = 2'b10;	 rom[1][30][5] = 2'b10;	 rom[1][31][5] = 2'b00;	 rom[1][32][5] = 2'b00;	 rom[1][33][5] = 2'b00;	 rom[1][34][5] = 2'b00;	 rom[1][35][5] = 2'b00;	 rom[1][36][5] = 2'b00;	 rom[1][37][5] = 2'b00;	 rom[1][38][5] = 2'b00;	 rom[1][39][5] = 2'b00;
 rom[1][0][6] = 2'b00;	 rom[1][1][6] = 2'b00;	 rom[1][2][6] = 2'b00;	 rom[1][3][6] = 2'b00;	 rom[1][4][6] = 2'b00;	 rom[1][5][6] = 2'b00;	 rom[1][6][6] = 2'b00;	 rom[1][7][6] = 2'b00;	 rom[1][8][6] = 2'b10;	 rom[1][9][6] = 2'b10;	 rom[1][10][6] = 2'b10;	 rom[1][11][6] = 2'b10;	 rom[1][12][6] = 2'b11;	 rom[1][13][6] = 2'b11;	 rom[1][14][6] = 2'b11;	 rom[1][15][6] = 2'b10;	 rom[1][16][6] = 2'b10;	 rom[1][17][6] = 2'b10;	 rom[1][18][6] = 2'b10;	 rom[1][19][6] = 2'b10;	 rom[1][20][6] = 2'b10;	 rom[1][21][6] = 2'b10;	 rom[1][22][6] = 2'b10;	 rom[1][23][6] = 2'b10;	 rom[1][24][6] = 2'b10;	 rom[1][25][6] = 2'b11;	 rom[1][26][6] = 2'b11;	 rom[1][27][6] = 2'b11;	 rom[1][28][6] = 2'b10;	 rom[1][29][6] = 2'b10;	 rom[1][30][6] = 2'b10;	 rom[1][31][6] = 2'b10;	 rom[1][32][6] = 2'b00;	 rom[1][33][6] = 2'b00;	 rom[1][34][6] = 2'b00;	 rom[1][35][6] = 2'b00;	 rom[1][36][6] = 2'b00;	 rom[1][37][6] = 2'b00;	 rom[1][38][6] = 2'b00;	 rom[1][39][6] = 2'b00;
 rom[1][0][7] = 2'b00;	 rom[1][1][7] = 2'b00;	 rom[1][2][7] = 2'b00;	 rom[1][3][7] = 2'b00;	 rom[1][4][7] = 2'b00;	 rom[1][5][7] = 2'b00;	 rom[1][6][7] = 2'b00;	 rom[1][7][7] = 2'b00;	 rom[1][8][7] = 2'b10;	 rom[1][9][7] = 2'b10;	 rom[1][10][7] = 2'b10;	 rom[1][11][7] = 2'b10;	 rom[1][12][7] = 2'b10;	 rom[1][13][7] = 2'b11;	 rom[1][14][7] = 2'b11;	 rom[1][15][7] = 2'b10;	 rom[1][16][7] = 2'b10;	 rom[1][17][7] = 2'b10;	 rom[1][18][7] = 2'b10;	 rom[1][19][7] = 2'b10;	 rom[1][20][7] = 2'b10;	 rom[1][21][7] = 2'b10;	 rom[1][22][7] = 2'b10;	 rom[1][23][7] = 2'b10;	 rom[1][24][7] = 2'b10;	 rom[1][25][7] = 2'b11;	 rom[1][26][7] = 2'b11;	 rom[1][27][7] = 2'b10;	 rom[1][28][7] = 2'b10;	 rom[1][29][7] = 2'b10;	 rom[1][30][7] = 2'b10;	 rom[1][31][7] = 2'b10;	 rom[1][32][7] = 2'b00;	 rom[1][33][7] = 2'b00;	 rom[1][34][7] = 2'b00;	 rom[1][35][7] = 2'b00;	 rom[1][36][7] = 2'b00;	 rom[1][37][7] = 2'b00;	 rom[1][38][7] = 2'b00;	 rom[1][39][7] = 2'b00;
 rom[1][0][8] = 2'b00;	 rom[1][1][8] = 2'b00;	 rom[1][2][8] = 2'b00;	 rom[1][3][8] = 2'b00;	 rom[1][4][8] = 2'b00;	 rom[1][5][8] = 2'b00;	 rom[1][6][8] = 2'b00;	 rom[1][7][8] = 2'b00;	 rom[1][8][8] = 2'b10;	 rom[1][9][8] = 2'b10;	 rom[1][10][8] = 2'b10;	 rom[1][11][8] = 2'b10;	 rom[1][12][8] = 2'b10;	 rom[1][13][8] = 2'b11;	 rom[1][14][8] = 2'b11;	 rom[1][15][8] = 2'b10;	 rom[1][16][8] = 2'b10;	 rom[1][17][8] = 2'b10;	 rom[1][18][8] = 2'b10;	 rom[1][19][8] = 2'b10;	 rom[1][20][8] = 2'b10;	 rom[1][21][8] = 2'b10;	 rom[1][22][8] = 2'b10;	 rom[1][23][8] = 2'b10;	 rom[1][24][8] = 2'b10;	 rom[1][25][8] = 2'b11;	 rom[1][26][8] = 2'b11;	 rom[1][27][8] = 2'b10;	 rom[1][28][8] = 2'b10;	 rom[1][29][8] = 2'b10;	 rom[1][30][8] = 2'b10;	 rom[1][31][8] = 2'b10;	 rom[1][32][8] = 2'b00;	 rom[1][33][8] = 2'b00;	 rom[1][34][8] = 2'b00;	 rom[1][35][8] = 2'b00;	 rom[1][36][8] = 2'b00;	 rom[1][37][8] = 2'b00;	 rom[1][38][8] = 2'b00;	 rom[1][39][8] = 2'b00;
 rom[1][0][9] = 2'b00;	 rom[1][1][9] = 2'b00;	 rom[1][2][9] = 2'b00;	 rom[1][3][9] = 2'b00;	 rom[1][4][9] = 2'b10;	 rom[1][5][9] = 2'b10;	 rom[1][6][9] = 2'b10;	 rom[1][7][9] = 2'b10;	 rom[1][8][9] = 2'b10;	 rom[1][9][9] = 2'b10;	 rom[1][10][9] = 2'b10;	 rom[1][11][9] = 2'b10;	 rom[1][12][9] = 2'b10;	 rom[1][13][9] = 2'b10;	 rom[1][14][9] = 2'b10;	 rom[1][15][9] = 2'b10;	 rom[1][16][9] = 2'b01;	 rom[1][17][9] = 2'b01;	 rom[1][18][9] = 2'b01;	 rom[1][19][9] = 2'b01;	 rom[1][20][9] = 2'b01;	 rom[1][21][9] = 2'b01;	 rom[1][22][9] = 2'b01;	 rom[1][23][9] = 2'b01;	 rom[1][24][9] = 2'b10;	 rom[1][25][9] = 2'b10;	 rom[1][26][9] = 2'b10;	 rom[1][27][9] = 2'b10;	 rom[1][28][9] = 2'b10;	 rom[1][29][9] = 2'b10;	 rom[1][30][9] = 2'b10;	 rom[1][31][9] = 2'b10;	 rom[1][32][9] = 2'b10;	 rom[1][33][9] = 2'b10;	 rom[1][34][9] = 2'b10;	 rom[1][35][9] = 2'b10;	 rom[1][36][9] = 2'b00;	 rom[1][37][9] = 2'b00;	 rom[1][38][9] = 2'b00;	 rom[1][39][9] = 2'b00;
 rom[1][0][10] = 2'b00;	 rom[1][1][10] = 2'b00;	 rom[1][2][10] = 2'b00;	 rom[1][3][10] = 2'b10;	 rom[1][4][10] = 2'b10;	 rom[1][5][10] = 2'b10;	 rom[1][6][10] = 2'b10;	 rom[1][7][10] = 2'b10;	 rom[1][8][10] = 2'b10;	 rom[1][9][10] = 2'b10;	 rom[1][10][10] = 2'b10;	 rom[1][11][10] = 2'b10;	 rom[1][12][10] = 2'b01;	 rom[1][13][10] = 2'b01;	 rom[1][14][10] = 2'b01;	 rom[1][15][10] = 2'b01;	 rom[1][16][10] = 2'b01;	 rom[1][17][10] = 2'b01;	 rom[1][18][10] = 2'b01;	 rom[1][19][10] = 2'b01;	 rom[1][20][10] = 2'b01;	 rom[1][21][10] = 2'b01;	 rom[1][22][10] = 2'b01;	 rom[1][23][10] = 2'b01;	 rom[1][24][10] = 2'b01;	 rom[1][25][10] = 2'b01;	 rom[1][26][10] = 2'b01;	 rom[1][27][10] = 2'b01;	 rom[1][28][10] = 2'b10;	 rom[1][29][10] = 2'b10;	 rom[1][30][10] = 2'b10;	 rom[1][31][10] = 2'b10;	 rom[1][32][10] = 2'b10;	 rom[1][33][10] = 2'b10;	 rom[1][34][10] = 2'b10;	 rom[1][35][10] = 2'b10;	 rom[1][36][10] = 2'b10;	 rom[1][37][10] = 2'b00;	 rom[1][38][10] = 2'b00;	 rom[1][39][10] = 2'b00;
 rom[1][0][11] = 2'b00;	 rom[1][1][11] = 2'b00;	 rom[1][2][11] = 2'b10;	 rom[1][3][11] = 2'b10;	 rom[1][4][11] = 2'b01;	 rom[1][5][11] = 2'b01;	 rom[1][6][11] = 2'b01;	 rom[1][7][11] = 2'b01;	 rom[1][8][11] = 2'b10;	 rom[1][9][11] = 2'b10;	 rom[1][10][11] = 2'b10;	 rom[1][11][11] = 2'b01;	 rom[1][12][11] = 2'b01;	 rom[1][13][11] = 2'b01;	 rom[1][14][11] = 2'b01;	 rom[1][15][11] = 2'b01;	 rom[1][16][11] = 2'b01;	 rom[1][17][11] = 2'b01;	 rom[1][18][11] = 2'b01;	 rom[1][19][11] = 2'b01;	 rom[1][20][11] = 2'b01;	 rom[1][21][11] = 2'b01;	 rom[1][22][11] = 2'b01;	 rom[1][23][11] = 2'b01;	 rom[1][24][11] = 2'b01;	 rom[1][25][11] = 2'b01;	 rom[1][26][11] = 2'b01;	 rom[1][27][11] = 2'b01;	 rom[1][28][11] = 2'b01;	 rom[1][29][11] = 2'b10;	 rom[1][30][11] = 2'b10;	 rom[1][31][11] = 2'b10;	 rom[1][32][11] = 2'b01;	 rom[1][33][11] = 2'b01;	 rom[1][34][11] = 2'b01;	 rom[1][35][11] = 2'b01;	 rom[1][36][11] = 2'b10;	 rom[1][37][11] = 2'b10;	 rom[1][38][11] = 2'b00;	 rom[1][39][11] = 2'b00;
 rom[1][0][12] = 2'b00;	 rom[1][1][12] = 2'b00;	 rom[1][2][12] = 2'b10;	 rom[1][3][12] = 2'b01;	 rom[1][4][12] = 2'b01;	 rom[1][5][12] = 2'b01;	 rom[1][6][12] = 2'b01;	 rom[1][7][12] = 2'b10;	 rom[1][8][12] = 2'b10;	 rom[1][9][12] = 2'b10;	 rom[1][10][12] = 2'b01;	 rom[1][11][12] = 2'b01;	 rom[1][12][12] = 2'b01;	 rom[1][13][12] = 2'b01;	 rom[1][14][12] = 2'b01;	 rom[1][15][12] = 2'b01;	 rom[1][16][12] = 2'b01;	 rom[1][17][12] = 2'b01;	 rom[1][18][12] = 2'b01;	 rom[1][19][12] = 2'b01;	 rom[1][20][12] = 2'b01;	 rom[1][21][12] = 2'b01;	 rom[1][22][12] = 2'b01;	 rom[1][23][12] = 2'b01;	 rom[1][24][12] = 2'b01;	 rom[1][25][12] = 2'b01;	 rom[1][26][12] = 2'b01;	 rom[1][27][12] = 2'b01;	 rom[1][28][12] = 2'b01;	 rom[1][29][12] = 2'b01;	 rom[1][30][12] = 2'b10;	 rom[1][31][12] = 2'b10;	 rom[1][32][12] = 2'b10;	 rom[1][33][12] = 2'b01;	 rom[1][34][12] = 2'b01;	 rom[1][35][12] = 2'b01;	 rom[1][36][12] = 2'b01;	 rom[1][37][12] = 2'b10;	 rom[1][38][12] = 2'b00;	 rom[1][39][12] = 2'b00;
 rom[1][0][13] = 2'b00;	 rom[1][1][13] = 2'b00;	 rom[1][2][13] = 2'b10;	 rom[1][3][13] = 2'b01;	 rom[1][4][13] = 2'b01;	 rom[1][5][13] = 2'b01;	 rom[1][6][13] = 2'b10;	 rom[1][7][13] = 2'b10;	 rom[1][8][13] = 2'b10;	 rom[1][9][13] = 2'b01;	 rom[1][10][13] = 2'b01;	 rom[1][11][13] = 2'b01;	 rom[1][12][13] = 2'b01;	 rom[1][13][13] = 2'b01;	 rom[1][14][13] = 2'b01;	 rom[1][15][13] = 2'b01;	 rom[1][16][13] = 2'b01;	 rom[1][17][13] = 2'b01;	 rom[1][18][13] = 2'b01;	 rom[1][19][13] = 2'b01;	 rom[1][20][13] = 2'b01;	 rom[1][21][13] = 2'b01;	 rom[1][22][13] = 2'b01;	 rom[1][23][13] = 2'b01;	 rom[1][24][13] = 2'b01;	 rom[1][25][13] = 2'b01;	 rom[1][26][13] = 2'b01;	 rom[1][27][13] = 2'b01;	 rom[1][28][13] = 2'b01;	 rom[1][29][13] = 2'b01;	 rom[1][30][13] = 2'b01;	 rom[1][31][13] = 2'b10;	 rom[1][32][13] = 2'b10;	 rom[1][33][13] = 2'b10;	 rom[1][34][13] = 2'b01;	 rom[1][35][13] = 2'b01;	 rom[1][36][13] = 2'b01;	 rom[1][37][13] = 2'b10;	 rom[1][38][13] = 2'b00;	 rom[1][39][13] = 2'b00;
 rom[1][0][14] = 2'b00;	 rom[1][1][14] = 2'b00;	 rom[1][2][14] = 2'b10;	 rom[1][3][14] = 2'b01;	 rom[1][4][14] = 2'b01;	 rom[1][5][14] = 2'b01;	 rom[1][6][14] = 2'b10;	 rom[1][7][14] = 2'b10;	 rom[1][8][14] = 2'b10;	 rom[1][9][14] = 2'b01;	 rom[1][10][14] = 2'b01;	 rom[1][11][14] = 2'b01;	 rom[1][12][14] = 2'b01;	 rom[1][13][14] = 2'b01;	 rom[1][14][14] = 2'b01;	 rom[1][15][14] = 2'b01;	 rom[1][16][14] = 2'b01;	 rom[1][17][14] = 2'b01;	 rom[1][18][14] = 2'b01;	 rom[1][19][14] = 2'b01;	 rom[1][20][14] = 2'b01;	 rom[1][21][14] = 2'b01;	 rom[1][22][14] = 2'b01;	 rom[1][23][14] = 2'b01;	 rom[1][24][14] = 2'b01;	 rom[1][25][14] = 2'b01;	 rom[1][26][14] = 2'b01;	 rom[1][27][14] = 2'b01;	 rom[1][28][14] = 2'b01;	 rom[1][29][14] = 2'b01;	 rom[1][30][14] = 2'b01;	 rom[1][31][14] = 2'b01;	 rom[1][32][14] = 2'b10;	 rom[1][33][14] = 2'b10;	 rom[1][34][14] = 2'b01;	 rom[1][35][14] = 2'b01;	 rom[1][36][14] = 2'b01;	 rom[1][37][14] = 2'b10;	 rom[1][38][14] = 2'b00;	 rom[1][39][14] = 2'b00;
 rom[1][0][15] = 2'b00;	 rom[1][1][15] = 2'b00;	 rom[1][2][15] = 2'b10;	 rom[1][3][15] = 2'b01;	 rom[1][4][15] = 2'b01;	 rom[1][5][15] = 2'b01;	 rom[1][6][15] = 2'b10;	 rom[1][7][15] = 2'b10;	 rom[1][8][15] = 2'b01;	 rom[1][9][15] = 2'b01;	 rom[1][10][15] = 2'b01;	 rom[1][11][15] = 2'b01;	 rom[1][12][15] = 2'b01;	 rom[1][13][15] = 2'b01;	 rom[1][14][15] = 2'b01;	 rom[1][15][15] = 2'b01;	 rom[1][16][15] = 2'b01;	 rom[1][17][15] = 2'b01;	 rom[1][18][15] = 2'b01;	 rom[1][19][15] = 2'b01;	 rom[1][20][15] = 2'b01;	 rom[1][21][15] = 2'b01;	 rom[1][22][15] = 2'b01;	 rom[1][23][15] = 2'b01;	 rom[1][24][15] = 2'b01;	 rom[1][25][15] = 2'b01;	 rom[1][26][15] = 2'b01;	 rom[1][27][15] = 2'b01;	 rom[1][28][15] = 2'b01;	 rom[1][29][15] = 2'b01;	 rom[1][30][15] = 2'b01;	 rom[1][31][15] = 2'b01;	 rom[1][32][15] = 2'b10;	 rom[1][33][15] = 2'b10;	 rom[1][34][15] = 2'b01;	 rom[1][35][15] = 2'b01;	 rom[1][36][15] = 2'b01;	 rom[1][37][15] = 2'b10;	 rom[1][38][15] = 2'b00;	 rom[1][39][15] = 2'b00;
 rom[1][0][16] = 2'b00;	 rom[1][1][16] = 2'b00;	 rom[1][2][16] = 2'b10;	 rom[1][3][16] = 2'b01;	 rom[1][4][16] = 2'b01;	 rom[1][5][16] = 2'b01;	 rom[1][6][16] = 2'b10;	 rom[1][7][16] = 2'b10;	 rom[1][8][16] = 2'b01;	 rom[1][9][16] = 2'b01;	 rom[1][10][16] = 2'b01;	 rom[1][11][16] = 2'b01;	 rom[1][12][16] = 2'b01;	 rom[1][13][16] = 2'b01;	 rom[1][14][16] = 2'b01;	 rom[1][15][16] = 2'b01;	 rom[1][16][16] = 2'b01;	 rom[1][17][16] = 2'b01;	 rom[1][18][16] = 2'b01;	 rom[1][19][16] = 2'b01;	 rom[1][20][16] = 2'b01;	 rom[1][21][16] = 2'b01;	 rom[1][22][16] = 2'b01;	 rom[1][23][16] = 2'b01;	 rom[1][24][16] = 2'b01;	 rom[1][25][16] = 2'b01;	 rom[1][26][16] = 2'b01;	 rom[1][27][16] = 2'b01;	 rom[1][28][16] = 2'b01;	 rom[1][29][16] = 2'b01;	 rom[1][30][16] = 2'b01;	 rom[1][31][16] = 2'b01;	 rom[1][32][16] = 2'b10;	 rom[1][33][16] = 2'b10;	 rom[1][34][16] = 2'b01;	 rom[1][35][16] = 2'b01;	 rom[1][36][16] = 2'b01;	 rom[1][37][16] = 2'b10;	 rom[1][38][16] = 2'b00;	 rom[1][39][16] = 2'b00;
 rom[1][0][17] = 2'b00;	 rom[1][1][17] = 2'b00;	 rom[1][2][17] = 2'b10;	 rom[1][3][17] = 2'b01;	 rom[1][4][17] = 2'b01;	 rom[1][5][17] = 2'b01;	 rom[1][6][17] = 2'b10;	 rom[1][7][17] = 2'b10;	 rom[1][8][17] = 2'b10;	 rom[1][9][17] = 2'b01;	 rom[1][10][17] = 2'b01;	 rom[1][11][17] = 2'b01;	 rom[1][12][17] = 2'b01;	 rom[1][13][17] = 2'b01;	 rom[1][14][17] = 2'b01;	 rom[1][15][17] = 2'b01;	 rom[1][16][17] = 2'b01;	 rom[1][17][17] = 2'b01;	 rom[1][18][17] = 2'b01;	 rom[1][19][17] = 2'b01;	 rom[1][20][17] = 2'b01;	 rom[1][21][17] = 2'b01;	 rom[1][22][17] = 2'b01;	 rom[1][23][17] = 2'b01;	 rom[1][24][17] = 2'b01;	 rom[1][25][17] = 2'b01;	 rom[1][26][17] = 2'b01;	 rom[1][27][17] = 2'b01;	 rom[1][28][17] = 2'b01;	 rom[1][29][17] = 2'b01;	 rom[1][30][17] = 2'b01;	 rom[1][31][17] = 2'b01;	 rom[1][32][17] = 2'b10;	 rom[1][33][17] = 2'b10;	 rom[1][34][17] = 2'b01;	 rom[1][35][17] = 2'b01;	 rom[1][36][17] = 2'b01;	 rom[1][37][17] = 2'b10;	 rom[1][38][17] = 2'b00;	 rom[1][39][17] = 2'b00;
 rom[1][0][18] = 2'b00;	 rom[1][1][18] = 2'b00;	 rom[1][2][18] = 2'b10;	 rom[1][3][18] = 2'b01;	 rom[1][4][18] = 2'b01;	 rom[1][5][18] = 2'b01;	 rom[1][6][18] = 2'b10;	 rom[1][7][18] = 2'b10;	 rom[1][8][18] = 2'b01;	 rom[1][9][18] = 2'b01;	 rom[1][10][18] = 2'b01;	 rom[1][11][18] = 2'b01;	 rom[1][12][18] = 2'b01;	 rom[1][13][18] = 2'b01;	 rom[1][14][18] = 2'b01;	 rom[1][15][18] = 2'b01;	 rom[1][16][18] = 2'b01;	 rom[1][17][18] = 2'b01;	 rom[1][18][18] = 2'b01;	 rom[1][19][18] = 2'b01;	 rom[1][20][18] = 2'b01;	 rom[1][21][18] = 2'b01;	 rom[1][22][18] = 2'b01;	 rom[1][23][18] = 2'b01;	 rom[1][24][18] = 2'b01;	 rom[1][25][18] = 2'b01;	 rom[1][26][18] = 2'b01;	 rom[1][27][18] = 2'b01;	 rom[1][28][18] = 2'b01;	 rom[1][29][18] = 2'b01;	 rom[1][30][18] = 2'b01;	 rom[1][31][18] = 2'b01;	 rom[1][32][18] = 2'b10;	 rom[1][33][18] = 2'b10;	 rom[1][34][18] = 2'b01;	 rom[1][35][18] = 2'b01;	 rom[1][36][18] = 2'b01;	 rom[1][37][18] = 2'b10;	 rom[1][38][18] = 2'b00;	 rom[1][39][18] = 2'b00;
 rom[1][0][19] = 2'b00;	 rom[1][1][19] = 2'b00;	 rom[1][2][19] = 2'b10;	 rom[1][3][19] = 2'b01;	 rom[1][4][19] = 2'b01;	 rom[1][5][19] = 2'b01;	 rom[1][6][19] = 2'b10;	 rom[1][7][19] = 2'b10;	 rom[1][8][19] = 2'b01;	 rom[1][9][19] = 2'b01;	 rom[1][10][19] = 2'b01;	 rom[1][11][19] = 2'b01;	 rom[1][12][19] = 2'b01;	 rom[1][13][19] = 2'b01;	 rom[1][14][19] = 2'b01;	 rom[1][15][19] = 2'b01;	 rom[1][16][19] = 2'b01;	 rom[1][17][19] = 2'b01;	 rom[1][18][19] = 2'b01;	 rom[1][19][19] = 2'b01;	 rom[1][20][19] = 2'b01;	 rom[1][21][19] = 2'b01;	 rom[1][22][19] = 2'b01;	 rom[1][23][19] = 2'b01;	 rom[1][24][19] = 2'b01;	 rom[1][25][19] = 2'b01;	 rom[1][26][19] = 2'b01;	 rom[1][27][19] = 2'b01;	 rom[1][28][19] = 2'b01;	 rom[1][29][19] = 2'b01;	 rom[1][30][19] = 2'b01;	 rom[1][31][19] = 2'b01;	 rom[1][32][19] = 2'b10;	 rom[1][33][19] = 2'b10;	 rom[1][34][19] = 2'b01;	 rom[1][35][19] = 2'b01;	 rom[1][36][19] = 2'b10;	 rom[1][37][19] = 2'b10;	 rom[1][38][19] = 2'b00;	 rom[1][39][19] = 2'b00;
 rom[1][0][20] = 2'b00;	 rom[1][1][20] = 2'b00;	 rom[1][2][20] = 2'b10;	 rom[1][3][20] = 2'b01;	 rom[1][4][20] = 2'b01;	 rom[1][5][20] = 2'b01;	 rom[1][6][20] = 2'b10;	 rom[1][7][20] = 2'b10;	 rom[1][8][20] = 2'b10;	 rom[1][9][20] = 2'b01;	 rom[1][10][20] = 2'b01;	 rom[1][11][20] = 2'b01;	 rom[1][12][20] = 2'b01;	 rom[1][13][20] = 2'b01;	 rom[1][14][20] = 2'b01;	 rom[1][15][20] = 2'b01;	 rom[1][16][20] = 2'b01;	 rom[1][17][20] = 2'b01;	 rom[1][18][20] = 2'b01;	 rom[1][19][20] = 2'b01;	 rom[1][20][20] = 2'b01;	 rom[1][21][20] = 2'b01;	 rom[1][22][20] = 2'b01;	 rom[1][23][20] = 2'b01;	 rom[1][24][20] = 2'b01;	 rom[1][25][20] = 2'b01;	 rom[1][26][20] = 2'b01;	 rom[1][27][20] = 2'b01;	 rom[1][28][20] = 2'b01;	 rom[1][29][20] = 2'b01;	 rom[1][30][20] = 2'b01;	 rom[1][31][20] = 2'b10;	 rom[1][32][20] = 2'b10;	 rom[1][33][20] = 2'b10;	 rom[1][34][20] = 2'b01;	 rom[1][35][20] = 2'b10;	 rom[1][36][20] = 2'b10;	 rom[1][37][20] = 2'b10;	 rom[1][38][20] = 2'b00;	 rom[1][39][20] = 2'b00;
 rom[1][0][21] = 2'b00;	 rom[1][1][21] = 2'b00;	 rom[1][2][21] = 2'b10;	 rom[1][3][21] = 2'b01;	 rom[1][4][21] = 2'b01;	 rom[1][5][21] = 2'b01;	 rom[1][6][21] = 2'b10;	 rom[1][7][21] = 2'b10;	 rom[1][8][21] = 2'b10;	 rom[1][9][21] = 2'b01;	 rom[1][10][21] = 2'b01;	 rom[1][11][21] = 2'b01;	 rom[1][12][21] = 2'b01;	 rom[1][13][21] = 2'b01;	 rom[1][14][21] = 2'b01;	 rom[1][15][21] = 2'b01;	 rom[1][16][21] = 2'b01;	 rom[1][17][21] = 2'b01;	 rom[1][18][21] = 2'b01;	 rom[1][19][21] = 2'b01;	 rom[1][20][21] = 2'b01;	 rom[1][21][21] = 2'b01;	 rom[1][22][21] = 2'b01;	 rom[1][23][21] = 2'b01;	 rom[1][24][21] = 2'b01;	 rom[1][25][21] = 2'b01;	 rom[1][26][21] = 2'b01;	 rom[1][27][21] = 2'b01;	 rom[1][28][21] = 2'b01;	 rom[1][29][21] = 2'b01;	 rom[1][30][21] = 2'b01;	 rom[1][31][21] = 2'b10;	 rom[1][32][21] = 2'b10;	 rom[1][33][21] = 2'b10;	 rom[1][34][21] = 2'b10;	 rom[1][35][21] = 2'b10;	 rom[1][36][21] = 2'b00;	 rom[1][37][21] = 2'b00;	 rom[1][38][21] = 2'b00;	 rom[1][39][21] = 2'b00;
 rom[1][0][22] = 2'b00;	 rom[1][1][22] = 2'b00;	 rom[1][2][22] = 2'b10;	 rom[1][3][22] = 2'b01;	 rom[1][4][22] = 2'b01;	 rom[1][5][22] = 2'b01;	 rom[1][6][22] = 2'b10;	 rom[1][7][22] = 2'b10;	 rom[1][8][22] = 2'b10;	 rom[1][9][22] = 2'b01;	 rom[1][10][22] = 2'b01;	 rom[1][11][22] = 2'b01;	 rom[1][12][22] = 2'b01;	 rom[1][13][22] = 2'b01;	 rom[1][14][22] = 2'b01;	 rom[1][15][22] = 2'b01;	 rom[1][16][22] = 2'b01;	 rom[1][17][22] = 2'b01;	 rom[1][18][22] = 2'b01;	 rom[1][19][22] = 2'b01;	 rom[1][20][22] = 2'b01;	 rom[1][21][22] = 2'b01;	 rom[1][22][22] = 2'b01;	 rom[1][23][22] = 2'b01;	 rom[1][24][22] = 2'b01;	 rom[1][25][22] = 2'b01;	 rom[1][26][22] = 2'b01;	 rom[1][27][22] = 2'b01;	 rom[1][28][22] = 2'b01;	 rom[1][29][22] = 2'b01;	 rom[1][30][22] = 2'b01;	 rom[1][31][22] = 2'b10;	 rom[1][32][22] = 2'b10;	 rom[1][33][22] = 2'b10;	 rom[1][34][22] = 2'b00;	 rom[1][35][22] = 2'b00;	 rom[1][36][22] = 2'b00;	 rom[1][37][22] = 2'b00;	 rom[1][38][22] = 2'b00;	 rom[1][39][22] = 2'b00;
 rom[1][0][23] = 2'b00;	 rom[1][1][23] = 2'b00;	 rom[1][2][23] = 2'b10;	 rom[1][3][23] = 2'b01;	 rom[1][4][23] = 2'b01;	 rom[1][5][23] = 2'b01;	 rom[1][6][23] = 2'b10;	 rom[1][7][23] = 2'b10;	 rom[1][8][23] = 2'b10;	 rom[1][9][23] = 2'b10;	 rom[1][10][23] = 2'b01;	 rom[1][11][23] = 2'b01;	 rom[1][12][23] = 2'b01;	 rom[1][13][23] = 2'b01;	 rom[1][14][23] = 2'b01;	 rom[1][15][23] = 2'b01;	 rom[1][16][23] = 2'b01;	 rom[1][17][23] = 2'b01;	 rom[1][18][23] = 2'b01;	 rom[1][19][23] = 2'b01;	 rom[1][20][23] = 2'b01;	 rom[1][21][23] = 2'b01;	 rom[1][22][23] = 2'b01;	 rom[1][23][23] = 2'b01;	 rom[1][24][23] = 2'b01;	 rom[1][25][23] = 2'b01;	 rom[1][26][23] = 2'b01;	 rom[1][27][23] = 2'b01;	 rom[1][28][23] = 2'b01;	 rom[1][29][23] = 2'b01;	 rom[1][30][23] = 2'b10;	 rom[1][31][23] = 2'b10;	 rom[1][32][23] = 2'b00;	 rom[1][33][23] = 2'b00;	 rom[1][34][23] = 2'b00;	 rom[1][35][23] = 2'b00;	 rom[1][36][23] = 2'b00;	 rom[1][37][23] = 2'b00;	 rom[1][38][23] = 2'b00;	 rom[1][39][23] = 2'b00;
 rom[1][0][24] = 2'b10;	 rom[1][1][24] = 2'b10;	 rom[1][2][24] = 2'b10;	 rom[1][3][24] = 2'b01;	 rom[1][4][24] = 2'b01;	 rom[1][5][24] = 2'b01;	 rom[1][6][24] = 2'b10;	 rom[1][7][24] = 2'b10;	 rom[1][8][24] = 2'b11;	 rom[1][9][24] = 2'b10;	 rom[1][10][24] = 2'b10;	 rom[1][11][24] = 2'b01;	 rom[1][12][24] = 2'b01;	 rom[1][13][24] = 2'b01;	 rom[1][14][24] = 2'b01;	 rom[1][15][24] = 2'b01;	 rom[1][16][24] = 2'b01;	 rom[1][17][24] = 2'b01;	 rom[1][18][24] = 2'b01;	 rom[1][19][24] = 2'b01;	 rom[1][20][24] = 2'b01;	 rom[1][21][24] = 2'b01;	 rom[1][22][24] = 2'b01;	 rom[1][23][24] = 2'b01;	 rom[1][24][24] = 2'b01;	 rom[1][25][24] = 2'b01;	 rom[1][26][24] = 2'b01;	 rom[1][27][24] = 2'b01;	 rom[1][28][24] = 2'b01;	 rom[1][29][24] = 2'b10;	 rom[1][30][24] = 2'b10;	 rom[1][31][24] = 2'b10;	 rom[1][32][24] = 2'b10;	 rom[1][33][24] = 2'b00;	 rom[1][34][24] = 2'b00;	 rom[1][35][24] = 2'b00;	 rom[1][36][24] = 2'b00;	 rom[1][37][24] = 2'b00;	 rom[1][38][24] = 2'b00;	 rom[1][39][24] = 2'b00;
 rom[1][0][25] = 2'b10;	 rom[1][1][25] = 2'b11;	 rom[1][2][25] = 2'b10;	 rom[1][3][25] = 2'b10;	 rom[1][4][25] = 2'b01;	 rom[1][5][25] = 2'b01;	 rom[1][6][25] = 2'b10;	 rom[1][7][25] = 2'b10;	 rom[1][8][25] = 2'b11;	 rom[1][9][25] = 2'b11;	 rom[1][10][25] = 2'b10;	 rom[1][11][25] = 2'b10;	 rom[1][12][25] = 2'b01;	 rom[1][13][25] = 2'b01;	 rom[1][14][25] = 2'b01;	 rom[1][15][25] = 2'b01;	 rom[1][16][25] = 2'b01;	 rom[1][17][25] = 2'b01;	 rom[1][18][25] = 2'b01;	 rom[1][19][25] = 2'b01;	 rom[1][20][25] = 2'b01;	 rom[1][21][25] = 2'b01;	 rom[1][22][25] = 2'b01;	 rom[1][23][25] = 2'b01;	 rom[1][24][25] = 2'b01;	 rom[1][25][25] = 2'b01;	 rom[1][26][25] = 2'b01;	 rom[1][27][25] = 2'b01;	 rom[1][28][25] = 2'b10;	 rom[1][29][25] = 2'b10;	 rom[1][30][25] = 2'b10;	 rom[1][31][25] = 2'b11;	 rom[1][32][25] = 2'b10;	 rom[1][33][25] = 2'b00;	 rom[1][34][25] = 2'b00;	 rom[1][35][25] = 2'b00;	 rom[1][36][25] = 2'b00;	 rom[1][37][25] = 2'b00;	 rom[1][38][25] = 2'b00;	 rom[1][39][25] = 2'b00;
 rom[1][0][26] = 2'b10;	 rom[1][1][26] = 2'b11;	 rom[1][2][26] = 2'b11;	 rom[1][3][26] = 2'b10;	 rom[1][4][26] = 2'b01;	 rom[1][5][26] = 2'b01;	 rom[1][6][26] = 2'b01;	 rom[1][7][26] = 2'b10;	 rom[1][8][26] = 2'b11;	 rom[1][9][26] = 2'b11;	 rom[1][10][26] = 2'b10;	 rom[1][11][26] = 2'b10;	 rom[1][12][26] = 2'b10;	 rom[1][13][26] = 2'b01;	 rom[1][14][26] = 2'b01;	 rom[1][15][26] = 2'b01;	 rom[1][16][26] = 2'b01;	 rom[1][17][26] = 2'b01;	 rom[1][18][26] = 2'b01;	 rom[1][19][26] = 2'b01;	 rom[1][20][26] = 2'b01;	 rom[1][21][26] = 2'b01;	 rom[1][22][26] = 2'b01;	 rom[1][23][26] = 2'b01;	 rom[1][24][26] = 2'b01;	 rom[1][25][26] = 2'b01;	 rom[1][26][26] = 2'b01;	 rom[1][27][26] = 2'b10;	 rom[1][28][26] = 2'b10;	 rom[1][29][26] = 2'b10;	 rom[1][30][26] = 2'b11;	 rom[1][31][26] = 2'b11;	 rom[1][32][26] = 2'b10;	 rom[1][33][26] = 2'b00;	 rom[1][34][26] = 2'b00;	 rom[1][35][26] = 2'b00;	 rom[1][36][26] = 2'b00;	 rom[1][37][26] = 2'b00;	 rom[1][38][26] = 2'b00;	 rom[1][39][26] = 2'b00;
 rom[1][0][27] = 2'b10;	 rom[1][1][27] = 2'b11;	 rom[1][2][27] = 2'b11;	 rom[1][3][27] = 2'b10;	 rom[1][4][27] = 2'b10;	 rom[1][5][27] = 2'b01;	 rom[1][6][27] = 2'b01;	 rom[1][7][27] = 2'b10;	 rom[1][8][27] = 2'b11;	 rom[1][9][27] = 2'b11;	 rom[1][10][27] = 2'b10;	 rom[1][11][27] = 2'b00;	 rom[1][12][27] = 2'b10;	 rom[1][13][27] = 2'b10;	 rom[1][14][27] = 2'b01;	 rom[1][15][27] = 2'b01;	 rom[1][16][27] = 2'b01;	 rom[1][17][27] = 2'b01;	 rom[1][18][27] = 2'b01;	 rom[1][19][27] = 2'b01;	 rom[1][20][27] = 2'b01;	 rom[1][21][27] = 2'b01;	 rom[1][22][27] = 2'b01;	 rom[1][23][27] = 2'b01;	 rom[1][24][27] = 2'b01;	 rom[1][25][27] = 2'b01;	 rom[1][26][27] = 2'b10;	 rom[1][27][27] = 2'b10;	 rom[1][28][27] = 2'b11;	 rom[1][29][27] = 2'b11;	 rom[1][30][27] = 2'b11;	 rom[1][31][27] = 2'b11;	 rom[1][32][27] = 2'b10;	 rom[1][33][27] = 2'b00;	 rom[1][34][27] = 2'b00;	 rom[1][35][27] = 2'b00;	 rom[1][36][27] = 2'b00;	 rom[1][37][27] = 2'b00;	 rom[1][38][27] = 2'b00;	 rom[1][39][27] = 2'b00;
 rom[1][0][28] = 2'b10;	 rom[1][1][28] = 2'b10;	 rom[1][2][28] = 2'b10;	 rom[1][3][28] = 2'b10;	 rom[1][4][28] = 2'b10;	 rom[1][5][28] = 2'b10;	 rom[1][6][28] = 2'b01;	 rom[1][7][28] = 2'b10;	 rom[1][8][28] = 2'b11;	 rom[1][9][28] = 2'b11;	 rom[1][10][28] = 2'b10;	 rom[1][11][28] = 2'b00;	 rom[1][12][28] = 2'b10;	 rom[1][13][28] = 2'b10;	 rom[1][14][28] = 2'b10;	 rom[1][15][28] = 2'b10;	 rom[1][16][28] = 2'b10;	 rom[1][17][28] = 2'b10;	 rom[1][18][28] = 2'b10;	 rom[1][19][28] = 2'b10;	 rom[1][20][28] = 2'b10;	 rom[1][21][28] = 2'b10;	 rom[1][22][28] = 2'b10;	 rom[1][23][28] = 2'b10;	 rom[1][24][28] = 2'b10;	 rom[1][25][28] = 2'b10;	 rom[1][26][28] = 2'b10;	 rom[1][27][28] = 2'b10;	 rom[1][28][28] = 2'b11;	 rom[1][29][28] = 2'b11;	 rom[1][30][28] = 2'b11;	 rom[1][31][28] = 2'b11;	 rom[1][32][28] = 2'b10;	 rom[1][33][28] = 2'b00;	 rom[1][34][28] = 2'b00;	 rom[1][35][28] = 2'b00;	 rom[1][36][28] = 2'b00;	 rom[1][37][28] = 2'b00;	 rom[1][38][28] = 2'b00;	 rom[1][39][28] = 2'b00;
 rom[1][0][29] = 2'b00;	 rom[1][1][29] = 2'b00;	 rom[1][2][29] = 2'b00;	 rom[1][3][29] = 2'b00;	 rom[1][4][29] = 2'b00;	 rom[1][5][29] = 2'b10;	 rom[1][6][29] = 2'b01;	 rom[1][7][29] = 2'b10;	 rom[1][8][29] = 2'b11;	 rom[1][9][29] = 2'b11;	 rom[1][10][29] = 2'b10;	 rom[1][11][29] = 2'b00;	 rom[1][12][29] = 2'b00;	 rom[1][13][29] = 2'b10;	 rom[1][14][29] = 2'b10;	 rom[1][15][29] = 2'b10;	 rom[1][16][29] = 2'b10;	 rom[1][17][29] = 2'b10;	 rom[1][18][29] = 2'b10;	 rom[1][19][29] = 2'b10;	 rom[1][20][29] = 2'b10;	 rom[1][21][29] = 2'b10;	 rom[1][22][29] = 2'b10;	 rom[1][23][29] = 2'b10;	 rom[1][24][29] = 2'b10;	 rom[1][25][29] = 2'b10;	 rom[1][26][29] = 2'b11;	 rom[1][27][29] = 2'b11;	 rom[1][28][29] = 2'b11;	 rom[1][29][29] = 2'b11;	 rom[1][30][29] = 2'b11;	 rom[1][31][29] = 2'b11;	 rom[1][32][29] = 2'b10;	 rom[1][33][29] = 2'b00;	 rom[1][34][29] = 2'b00;	 rom[1][35][29] = 2'b00;	 rom[1][36][29] = 2'b00;	 rom[1][37][29] = 2'b00;	 rom[1][38][29] = 2'b00;	 rom[1][39][29] = 2'b00;
 rom[1][0][30] = 2'b00;	 rom[1][1][30] = 2'b00;	 rom[1][2][30] = 2'b00;	 rom[1][3][30] = 2'b00;	 rom[1][4][30] = 2'b00;	 rom[1][5][30] = 2'b10;	 rom[1][6][30] = 2'b10;	 rom[1][7][30] = 2'b10;	 rom[1][8][30] = 2'b11;	 rom[1][9][30] = 2'b11;	 rom[1][10][30] = 2'b10;	 rom[1][11][30] = 2'b00;	 rom[1][12][30] = 2'b00;	 rom[1][13][30] = 2'b10;	 rom[1][14][30] = 2'b11;	 rom[1][15][30] = 2'b11;	 rom[1][16][30] = 2'b11;	 rom[1][17][30] = 2'b11;	 rom[1][18][30] = 2'b11;	 rom[1][19][30] = 2'b11;	 rom[1][20][30] = 2'b11;	 rom[1][21][30] = 2'b10;	 rom[1][22][30] = 2'b00;	 rom[1][23][30] = 2'b10;	 rom[1][24][30] = 2'b10;	 rom[1][25][30] = 2'b11;	 rom[1][26][30] = 2'b11;	 rom[1][27][30] = 2'b11;	 rom[1][28][30] = 2'b11;	 rom[1][29][30] = 2'b11;	 rom[1][30][30] = 2'b11;	 rom[1][31][30] = 2'b10;	 rom[1][32][30] = 2'b10;	 rom[1][33][30] = 2'b00;	 rom[1][34][30] = 2'b00;	 rom[1][35][30] = 2'b00;	 rom[1][36][30] = 2'b00;	 rom[1][37][30] = 2'b00;	 rom[1][38][30] = 2'b00;	 rom[1][39][30] = 2'b00;
 rom[1][0][31] = 2'b00;	 rom[1][1][31] = 2'b00;	 rom[1][2][31] = 2'b00;	 rom[1][3][31] = 2'b00;	 rom[1][4][31] = 2'b00;	 rom[1][5][31] = 2'b00;	 rom[1][6][31] = 2'b10;	 rom[1][7][31] = 2'b10;	 rom[1][8][31] = 2'b11;	 rom[1][9][31] = 2'b11;	 rom[1][10][31] = 2'b10;	 rom[1][11][31] = 2'b00;	 rom[1][12][31] = 2'b00;	 rom[1][13][31] = 2'b10;	 rom[1][14][31] = 2'b10;	 rom[1][15][31] = 2'b11;	 rom[1][16][31] = 2'b11;	 rom[1][17][31] = 2'b11;	 rom[1][18][31] = 2'b11;	 rom[1][19][31] = 2'b11;	 rom[1][20][31] = 2'b11;	 rom[1][21][31] = 2'b10;	 rom[1][22][31] = 2'b00;	 rom[1][23][31] = 2'b00;	 rom[1][24][31] = 2'b10;	 rom[1][25][31] = 2'b10;	 rom[1][26][31] = 2'b11;	 rom[1][27][31] = 2'b11;	 rom[1][28][31] = 2'b11;	 rom[1][29][31] = 2'b11;	 rom[1][30][31] = 2'b10;	 rom[1][31][31] = 2'b10;	 rom[1][32][31] = 2'b00;	 rom[1][33][31] = 2'b00;	 rom[1][34][31] = 2'b00;	 rom[1][35][31] = 2'b00;	 rom[1][36][31] = 2'b00;	 rom[1][37][31] = 2'b00;	 rom[1][38][31] = 2'b00;	 rom[1][39][31] = 2'b00;
 rom[1][0][32] = 2'b00;	 rom[1][1][32] = 2'b00;	 rom[1][2][32] = 2'b00;	 rom[1][3][32] = 2'b00;	 rom[1][4][32] = 2'b00;	 rom[1][5][32] = 2'b00;	 rom[1][6][32] = 2'b00;	 rom[1][7][32] = 2'b10;	 rom[1][8][32] = 2'b11;	 rom[1][9][32] = 2'b11;	 rom[1][10][32] = 2'b10;	 rom[1][11][32] = 2'b00;	 rom[1][12][32] = 2'b00;	 rom[1][13][32] = 2'b00;	 rom[1][14][32] = 2'b10;	 rom[1][15][32] = 2'b10;	 rom[1][16][32] = 2'b11;	 rom[1][17][32] = 2'b11;	 rom[1][18][32] = 2'b11;	 rom[1][19][32] = 2'b11;	 rom[1][20][32] = 2'b10;	 rom[1][21][32] = 2'b10;	 rom[1][22][32] = 2'b00;	 rom[1][23][32] = 2'b00;	 rom[1][24][32] = 2'b00;	 rom[1][25][32] = 2'b10;	 rom[1][26][32] = 2'b10;	 rom[1][27][32] = 2'b10;	 rom[1][28][32] = 2'b10;	 rom[1][29][32] = 2'b10;	 rom[1][30][32] = 2'b10;	 rom[1][31][32] = 2'b00;	 rom[1][32][32] = 2'b00;	 rom[1][33][32] = 2'b00;	 rom[1][34][32] = 2'b00;	 rom[1][35][32] = 2'b00;	 rom[1][36][32] = 2'b00;	 rom[1][37][32] = 2'b00;	 rom[1][38][32] = 2'b00;	 rom[1][39][32] = 2'b00;
 rom[1][0][33] = 2'b00;	 rom[1][1][33] = 2'b00;	 rom[1][2][33] = 2'b00;	 rom[1][3][33] = 2'b00;	 rom[1][4][33] = 2'b00;	 rom[1][5][33] = 2'b00;	 rom[1][6][33] = 2'b00;	 rom[1][7][33] = 2'b10;	 rom[1][8][33] = 2'b11;	 rom[1][9][33] = 2'b11;	 rom[1][10][33] = 2'b10;	 rom[1][11][33] = 2'b00;	 rom[1][12][33] = 2'b00;	 rom[1][13][33] = 2'b00;	 rom[1][14][33] = 2'b00;	 rom[1][15][33] = 2'b10;	 rom[1][16][33] = 2'b10;	 rom[1][17][33] = 2'b10;	 rom[1][18][33] = 2'b10;	 rom[1][19][33] = 2'b10;	 rom[1][20][33] = 2'b10;	 rom[1][21][33] = 2'b00;	 rom[1][22][33] = 2'b00;	 rom[1][23][33] = 2'b00;	 rom[1][24][33] = 2'b00;	 rom[1][25][33] = 2'b00;	 rom[1][26][33] = 2'b00;	 rom[1][27][33] = 2'b00;	 rom[1][28][33] = 2'b00;	 rom[1][29][33] = 2'b00;	 rom[1][30][33] = 2'b00;	 rom[1][31][33] = 2'b00;	 rom[1][32][33] = 2'b00;	 rom[1][33][33] = 2'b00;	 rom[1][34][33] = 2'b00;	 rom[1][35][33] = 2'b00;	 rom[1][36][33] = 2'b00;	 rom[1][37][33] = 2'b00;	 rom[1][38][33] = 2'b00;	 rom[1][39][33] = 2'b00;
 rom[1][0][34] = 2'b00;	 rom[1][1][34] = 2'b00;	 rom[1][2][34] = 2'b00;	 rom[1][3][34] = 2'b00;	 rom[1][4][34] = 2'b00;	 rom[1][5][34] = 2'b00;	 rom[1][6][34] = 2'b00;	 rom[1][7][34] = 2'b10;	 rom[1][8][34] = 2'b11;	 rom[1][9][34] = 2'b11;	 rom[1][10][34] = 2'b10;	 rom[1][11][34] = 2'b00;	 rom[1][12][34] = 2'b00;	 rom[1][13][34] = 2'b00;	 rom[1][14][34] = 2'b00;	 rom[1][15][34] = 2'b00;	 rom[1][16][34] = 2'b00;	 rom[1][17][34] = 2'b00;	 rom[1][18][34] = 2'b00;	 rom[1][19][34] = 2'b00;	 rom[1][20][34] = 2'b00;	 rom[1][21][34] = 2'b00;	 rom[1][22][34] = 2'b00;	 rom[1][23][34] = 2'b00;	 rom[1][24][34] = 2'b00;	 rom[1][25][34] = 2'b00;	 rom[1][26][34] = 2'b00;	 rom[1][27][34] = 2'b00;	 rom[1][28][34] = 2'b00;	 rom[1][29][34] = 2'b00;	 rom[1][30][34] = 2'b00;	 rom[1][31][34] = 2'b00;	 rom[1][32][34] = 2'b00;	 rom[1][33][34] = 2'b00;	 rom[1][34][34] = 2'b00;	 rom[1][35][34] = 2'b00;	 rom[1][36][34] = 2'b00;	 rom[1][37][34] = 2'b00;	 rom[1][38][34] = 2'b00;	 rom[1][39][34] = 2'b00;
 rom[1][0][35] = 2'b00;	 rom[1][1][35] = 2'b00;	 rom[1][2][35] = 2'b00;	 rom[1][3][35] = 2'b00;	 rom[1][4][35] = 2'b00;	 rom[1][5][35] = 2'b00;	 rom[1][6][35] = 2'b00;	 rom[1][7][35] = 2'b10;	 rom[1][8][35] = 2'b11;	 rom[1][9][35] = 2'b11;	 rom[1][10][35] = 2'b10;	 rom[1][11][35] = 2'b00;	 rom[1][12][35] = 2'b00;	 rom[1][13][35] = 2'b00;	 rom[1][14][35] = 2'b00;	 rom[1][15][35] = 2'b00;	 rom[1][16][35] = 2'b00;	 rom[1][17][35] = 2'b00;	 rom[1][18][35] = 2'b00;	 rom[1][19][35] = 2'b00;	 rom[1][20][35] = 2'b00;	 rom[1][21][35] = 2'b00;	 rom[1][22][35] = 2'b00;	 rom[1][23][35] = 2'b00;	 rom[1][24][35] = 2'b00;	 rom[1][25][35] = 2'b00;	 rom[1][26][35] = 2'b00;	 rom[1][27][35] = 2'b00;	 rom[1][28][35] = 2'b00;	 rom[1][29][35] = 2'b00;	 rom[1][30][35] = 2'b00;	 rom[1][31][35] = 2'b00;	 rom[1][32][35] = 2'b00;	 rom[1][33][35] = 2'b00;	 rom[1][34][35] = 2'b00;	 rom[1][35][35] = 2'b00;	 rom[1][36][35] = 2'b00;	 rom[1][37][35] = 2'b00;	 rom[1][38][35] = 2'b00;	 rom[1][39][35] = 2'b00;
 rom[1][0][36] = 2'b00;	 rom[1][1][36] = 2'b00;	 rom[1][2][36] = 2'b00;	 rom[1][3][36] = 2'b00;	 rom[1][4][36] = 2'b00;	 rom[1][5][36] = 2'b00;	 rom[1][6][36] = 2'b00;	 rom[1][7][36] = 2'b10;	 rom[1][8][36] = 2'b11;	 rom[1][9][36] = 2'b11;	 rom[1][10][36] = 2'b10;	 rom[1][11][36] = 2'b00;	 rom[1][12][36] = 2'b00;	 rom[1][13][36] = 2'b00;	 rom[1][14][36] = 2'b00;	 rom[1][15][36] = 2'b00;	 rom[1][16][36] = 2'b00;	 rom[1][17][36] = 2'b00;	 rom[1][18][36] = 2'b00;	 rom[1][19][36] = 2'b00;	 rom[1][20][36] = 2'b00;	 rom[1][21][36] = 2'b00;	 rom[1][22][36] = 2'b00;	 rom[1][23][36] = 2'b00;	 rom[1][24][36] = 2'b00;	 rom[1][25][36] = 2'b00;	 rom[1][26][36] = 2'b00;	 rom[1][27][36] = 2'b00;	 rom[1][28][36] = 2'b00;	 rom[1][29][36] = 2'b00;	 rom[1][30][36] = 2'b00;	 rom[1][31][36] = 2'b00;	 rom[1][32][36] = 2'b00;	 rom[1][33][36] = 2'b00;	 rom[1][34][36] = 2'b00;	 rom[1][35][36] = 2'b00;	 rom[1][36][36] = 2'b00;	 rom[1][37][36] = 2'b00;	 rom[1][38][36] = 2'b00;	 rom[1][39][36] = 2'b00;
 rom[1][0][37] = 2'b00;	 rom[1][1][37] = 2'b00;	 rom[1][2][37] = 2'b00;	 rom[1][3][37] = 2'b00;	 rom[1][4][37] = 2'b00;	 rom[1][5][37] = 2'b00;	 rom[1][6][37] = 2'b00;	 rom[1][7][37] = 2'b10;	 rom[1][8][37] = 2'b11;	 rom[1][9][37] = 2'b11;	 rom[1][10][37] = 2'b10;	 rom[1][11][37] = 2'b00;	 rom[1][12][37] = 2'b00;	 rom[1][13][37] = 2'b00;	 rom[1][14][37] = 2'b00;	 rom[1][15][37] = 2'b00;	 rom[1][16][37] = 2'b00;	 rom[1][17][37] = 2'b00;	 rom[1][18][37] = 2'b00;	 rom[1][19][37] = 2'b00;	 rom[1][20][37] = 2'b00;	 rom[1][21][37] = 2'b00;	 rom[1][22][37] = 2'b00;	 rom[1][23][37] = 2'b00;	 rom[1][24][37] = 2'b00;	 rom[1][25][37] = 2'b00;	 rom[1][26][37] = 2'b00;	 rom[1][27][37] = 2'b00;	 rom[1][28][37] = 2'b00;	 rom[1][29][37] = 2'b00;	 rom[1][30][37] = 2'b00;	 rom[1][31][37] = 2'b00;	 rom[1][32][37] = 2'b00;	 rom[1][33][37] = 2'b00;	 rom[1][34][37] = 2'b00;	 rom[1][35][37] = 2'b00;	 rom[1][36][37] = 2'b00;	 rom[1][37][37] = 2'b00;	 rom[1][38][37] = 2'b00;	 rom[1][39][37] = 2'b00;
 rom[1][0][38] = 2'b00;	 rom[1][1][38] = 2'b00;	 rom[1][2][38] = 2'b00;	 rom[1][3][38] = 2'b00;	 rom[1][4][38] = 2'b00;	 rom[1][5][38] = 2'b00;	 rom[1][6][38] = 2'b10;	 rom[1][7][38] = 2'b10;	 rom[1][8][38] = 2'b11;	 rom[1][9][38] = 2'b11;	 rom[1][10][38] = 2'b10;	 rom[1][11][38] = 2'b10;	 rom[1][12][38] = 2'b00;	 rom[1][13][38] = 2'b00;	 rom[1][14][38] = 2'b00;	 rom[1][15][38] = 2'b00;	 rom[1][16][38] = 2'b00;	 rom[1][17][38] = 2'b00;	 rom[1][18][38] = 2'b00;	 rom[1][19][38] = 2'b00;	 rom[1][20][38] = 2'b00;	 rom[1][21][38] = 2'b00;	 rom[1][22][38] = 2'b00;	 rom[1][23][38] = 2'b00;	 rom[1][24][38] = 2'b00;	 rom[1][25][38] = 2'b00;	 rom[1][26][38] = 2'b00;	 rom[1][27][38] = 2'b00;	 rom[1][28][38] = 2'b00;	 rom[1][29][38] = 2'b00;	 rom[1][30][38] = 2'b00;	 rom[1][31][38] = 2'b00;	 rom[1][32][38] = 2'b00;	 rom[1][33][38] = 2'b00;	 rom[1][34][38] = 2'b00;	 rom[1][35][38] = 2'b00;	 rom[1][36][38] = 2'b00;	 rom[1][37][38] = 2'b00;	 rom[1][38][38] = 2'b00;	 rom[1][39][38] = 2'b00;
 rom[1][0][39] = 2'b00;	 rom[1][1][39] = 2'b00;	 rom[1][2][39] = 2'b00;	 rom[1][3][39] = 2'b00;	 rom[1][4][39] = 2'b00;	 rom[1][5][39] = 2'b00;	 rom[1][6][39] = 2'b10;	 rom[1][7][39] = 2'b10;	 rom[1][8][39] = 2'b10;	 rom[1][9][39] = 2'b10;	 rom[1][10][39] = 2'b10;	 rom[1][11][39] = 2'b10;	 rom[1][12][39] = 2'b00;	 rom[1][13][39] = 2'b00;	 rom[1][14][39] = 2'b00;	 rom[1][15][39] = 2'b00;	 rom[1][16][39] = 2'b00;	 rom[1][17][39] = 2'b00;	 rom[1][18][39] = 2'b00;	 rom[1][19][39] = 2'b00;	 rom[1][20][39] = 2'b00;	 rom[1][21][39] = 2'b00;	 rom[1][22][39] = 2'b00;	 rom[1][23][39] = 2'b00;	 rom[1][24][39] = 2'b00;	 rom[1][25][39] = 2'b00;	 rom[1][26][39] = 2'b00;	 rom[1][27][39] = 2'b00;	 rom[1][28][39] = 2'b00;	 rom[1][29][39] = 2'b00;	 rom[1][30][39] = 2'b00;	 rom[1][31][39] = 2'b00;	 rom[1][32][39] = 2'b00;	 rom[1][33][39] = 2'b00;	 rom[1][34][39] = 2'b00;	 rom[1][35][39] = 2'b00;	 rom[1][36][39] = 2'b00;	 rom[1][37][39] = 2'b00;	 rom[1][38][39] = 2'b00;	 rom[1][39][39] = 2'b00;
//left
 rom[2][0][0] = 2'b00;	 rom[2][1][0] = 2'b00;	 rom[2][2][0] = 2'b00;	 rom[2][3][0] = 2'b00;	 rom[2][4][0] = 2'b00;	 rom[2][5][0] = 2'b00;	 rom[2][6][0] = 2'b00;	 rom[2][7][0] = 2'b00;	 rom[2][8][0] = 2'b00;	 rom[2][9][0] = 2'b00;	 rom[2][10][0] = 2'b00;	 rom[2][11][0] = 2'b10;	 rom[2][12][0] = 2'b10;	 rom[2][13][0] = 2'b10;	 rom[2][14][0] = 2'b10;	 rom[2][15][0] = 2'b10;	 rom[2][16][0] = 2'b00;	 rom[2][17][0] = 2'b00;	 rom[2][18][0] = 2'b00;	 rom[2][19][0] = 2'b00;	 rom[2][20][0] = 2'b00;	 rom[2][21][0] = 2'b00;	 rom[2][22][0] = 2'b00;	 rom[2][23][0] = 2'b00;	 rom[2][24][0] = 2'b00;	 rom[2][25][0] = 2'b00;	 rom[2][26][0] = 2'b00;	 rom[2][27][0] = 2'b00;	 rom[2][28][0] = 2'b00;	 rom[2][29][0] = 2'b00;	 rom[2][30][0] = 2'b00;	 rom[2][31][0] = 2'b00;	 rom[2][32][0] = 2'b00;	 rom[2][33][0] = 2'b00;	 rom[2][34][0] = 2'b00;	 rom[2][35][0] = 2'b00;	 rom[2][36][0] = 2'b00;	 rom[2][37][0] = 2'b00;	 rom[2][38][0] = 2'b00;	 rom[2][39][0] = 2'b00;
 rom[2][0][1] = 2'b00;	 rom[2][1][1] = 2'b00;	 rom[2][2][1] = 2'b00;	 rom[2][3][1] = 2'b00;	 rom[2][4][1] = 2'b00;	 rom[2][5][1] = 2'b00;	 rom[2][6][1] = 2'b00;	 rom[2][7][1] = 2'b00;	 rom[2][8][1] = 2'b00;	 rom[2][9][1] = 2'b00;	 rom[2][10][1] = 2'b00;	 rom[2][11][1] = 2'b10;	 rom[2][12][1] = 2'b11;	 rom[2][13][1] = 2'b11;	 rom[2][14][1] = 2'b11;	 rom[2][15][1] = 2'b10;	 rom[2][16][1] = 2'b00;	 rom[2][17][1] = 2'b00;	 rom[2][18][1] = 2'b00;	 rom[2][19][1] = 2'b00;	 rom[2][20][1] = 2'b00;	 rom[2][21][1] = 2'b00;	 rom[2][22][1] = 2'b00;	 rom[2][23][1] = 2'b00;	 rom[2][24][1] = 2'b00;	 rom[2][25][1] = 2'b00;	 rom[2][26][1] = 2'b00;	 rom[2][27][1] = 2'b00;	 rom[2][28][1] = 2'b00;	 rom[2][29][1] = 2'b00;	 rom[2][30][1] = 2'b00;	 rom[2][31][1] = 2'b00;	 rom[2][32][1] = 2'b00;	 rom[2][33][1] = 2'b00;	 rom[2][34][1] = 2'b00;	 rom[2][35][1] = 2'b00;	 rom[2][36][1] = 2'b00;	 rom[2][37][1] = 2'b00;	 rom[2][38][1] = 2'b00;	 rom[2][39][1] = 2'b00;
 rom[2][0][2] = 2'b00;	 rom[2][1][2] = 2'b00;	 rom[2][2][2] = 2'b00;	 rom[2][3][2] = 2'b00;	 rom[2][4][2] = 2'b00;	 rom[2][5][2] = 2'b00;	 rom[2][6][2] = 2'b00;	 rom[2][7][2] = 2'b00;	 rom[2][8][2] = 2'b00;	 rom[2][9][2] = 2'b00;	 rom[2][10][2] = 2'b00;	 rom[2][11][2] = 2'b10;	 rom[2][12][2] = 2'b11;	 rom[2][13][2] = 2'b11;	 rom[2][14][2] = 2'b10;	 rom[2][15][2] = 2'b10;	 rom[2][16][2] = 2'b10;	 rom[2][17][2] = 2'b10;	 rom[2][18][2] = 2'b10;	 rom[2][19][2] = 2'b10;	 rom[2][20][2] = 2'b10;	 rom[2][21][2] = 2'b10;	 rom[2][22][2] = 2'b10;	 rom[2][23][2] = 2'b10;	 rom[2][24][2] = 2'b10;	 rom[2][25][2] = 2'b10;	 rom[2][26][2] = 2'b10;	 rom[2][27][2] = 2'b10;	 rom[2][28][2] = 2'b10;	 rom[2][29][2] = 2'b00;	 rom[2][30][2] = 2'b00;	 rom[2][31][2] = 2'b00;	 rom[2][32][2] = 2'b00;	 rom[2][33][2] = 2'b00;	 rom[2][34][2] = 2'b00;	 rom[2][35][2] = 2'b00;	 rom[2][36][2] = 2'b00;	 rom[2][37][2] = 2'b00;	 rom[2][38][2] = 2'b00;	 rom[2][39][2] = 2'b00;
 rom[2][0][3] = 2'b00;	 rom[2][1][3] = 2'b00;	 rom[2][2][3] = 2'b00;	 rom[2][3][3] = 2'b00;	 rom[2][4][3] = 2'b00;	 rom[2][5][3] = 2'b00;	 rom[2][6][3] = 2'b00;	 rom[2][7][3] = 2'b00;	 rom[2][8][3] = 2'b00;	 rom[2][9][3] = 2'b00;	 rom[2][10][3] = 2'b00;	 rom[2][11][3] = 2'b10;	 rom[2][12][3] = 2'b10;	 rom[2][13][3] = 2'b10;	 rom[2][14][3] = 2'b10;	 rom[2][15][3] = 2'b01;	 rom[2][16][3] = 2'b01;	 rom[2][17][3] = 2'b01;	 rom[2][18][3] = 2'b01;	 rom[2][19][3] = 2'b01;	 rom[2][20][3] = 2'b01;	 rom[2][21][3] = 2'b01;	 rom[2][22][3] = 2'b01;	 rom[2][23][3] = 2'b01;	 rom[2][24][3] = 2'b01;	 rom[2][25][3] = 2'b01;	 rom[2][26][3] = 2'b01;	 rom[2][27][3] = 2'b01;	 rom[2][28][3] = 2'b10;	 rom[2][29][3] = 2'b10;	 rom[2][30][3] = 2'b00;	 rom[2][31][3] = 2'b00;	 rom[2][32][3] = 2'b00;	 rom[2][33][3] = 2'b00;	 rom[2][34][3] = 2'b00;	 rom[2][35][3] = 2'b00;	 rom[2][36][3] = 2'b00;	 rom[2][37][3] = 2'b00;	 rom[2][38][3] = 2'b00;	 rom[2][39][3] = 2'b00;
 rom[2][0][4] = 2'b00;	 rom[2][1][4] = 2'b00;	 rom[2][2][4] = 2'b00;	 rom[2][3][4] = 2'b00;	 rom[2][4][4] = 2'b00;	 rom[2][5][4] = 2'b00;	 rom[2][6][4] = 2'b00;	 rom[2][7][4] = 2'b00;	 rom[2][8][4] = 2'b00;	 rom[2][9][4] = 2'b00;	 rom[2][10][4] = 2'b00;	 rom[2][11][4] = 2'b10;	 rom[2][12][4] = 2'b10;	 rom[2][13][4] = 2'b01;	 rom[2][14][4] = 2'b01;	 rom[2][15][4] = 2'b01;	 rom[2][16][4] = 2'b01;	 rom[2][17][4] = 2'b01;	 rom[2][18][4] = 2'b01;	 rom[2][19][4] = 2'b01;	 rom[2][20][4] = 2'b01;	 rom[2][21][4] = 2'b01;	 rom[2][22][4] = 2'b01;	 rom[2][23][4] = 2'b01;	 rom[2][24][4] = 2'b01;	 rom[2][25][4] = 2'b01;	 rom[2][26][4] = 2'b01;	 rom[2][27][4] = 2'b01;	 rom[2][28][4] = 2'b01;	 rom[2][29][4] = 2'b10;	 rom[2][30][4] = 2'b10;	 rom[2][31][4] = 2'b00;	 rom[2][32][4] = 2'b00;	 rom[2][33][4] = 2'b00;	 rom[2][34][4] = 2'b00;	 rom[2][35][4] = 2'b00;	 rom[2][36][4] = 2'b00;	 rom[2][37][4] = 2'b00;	 rom[2][38][4] = 2'b00;	 rom[2][39][4] = 2'b00;
 rom[2][0][5] = 2'b00;	 rom[2][1][5] = 2'b00;	 rom[2][2][5] = 2'b00;	 rom[2][3][5] = 2'b00;	 rom[2][4][5] = 2'b00;	 rom[2][5][5] = 2'b00;	 rom[2][6][5] = 2'b00;	 rom[2][7][5] = 2'b00;	 rom[2][8][5] = 2'b00;	 rom[2][9][5] = 2'b10;	 rom[2][10][5] = 2'b10;	 rom[2][11][5] = 2'b10;	 rom[2][12][5] = 2'b01;	 rom[2][13][5] = 2'b01;	 rom[2][14][5] = 2'b01;	 rom[2][15][5] = 2'b01;	 rom[2][16][5] = 2'b01;	 rom[2][17][5] = 2'b01;	 rom[2][18][5] = 2'b01;	 rom[2][19][5] = 2'b01;	 rom[2][20][5] = 2'b01;	 rom[2][21][5] = 2'b01;	 rom[2][22][5] = 2'b01;	 rom[2][23][5] = 2'b01;	 rom[2][24][5] = 2'b01;	 rom[2][25][5] = 2'b01;	 rom[2][26][5] = 2'b01;	 rom[2][27][5] = 2'b01;	 rom[2][28][5] = 2'b01;	 rom[2][29][5] = 2'b10;	 rom[2][30][5] = 2'b10;	 rom[2][31][5] = 2'b00;	 rom[2][32][5] = 2'b00;	 rom[2][33][5] = 2'b00;	 rom[2][34][5] = 2'b00;	 rom[2][35][5] = 2'b00;	 rom[2][36][5] = 2'b00;	 rom[2][37][5] = 2'b00;	 rom[2][38][5] = 2'b00;	 rom[2][39][5] = 2'b00;
 rom[2][0][6] = 2'b10;	 rom[2][1][6] = 2'b10;	 rom[2][2][6] = 2'b00;	 rom[2][3][6] = 2'b00;	 rom[2][4][6] = 2'b00;	 rom[2][5][6] = 2'b00;	 rom[2][6][6] = 2'b00;	 rom[2][7][6] = 2'b00;	 rom[2][8][6] = 2'b10;	 rom[2][9][6] = 2'b10;	 rom[2][10][6] = 2'b01;	 rom[2][11][6] = 2'b01;	 rom[2][12][6] = 2'b01;	 rom[2][13][6] = 2'b01;	 rom[2][14][6] = 2'b10;	 rom[2][15][6] = 2'b10;	 rom[2][16][6] = 2'b10;	 rom[2][17][6] = 2'b10;	 rom[2][18][6] = 2'b10;	 rom[2][19][6] = 2'b10;	 rom[2][20][6] = 2'b10;	 rom[2][21][6] = 2'b10;	 rom[2][22][6] = 2'b10;	 rom[2][23][6] = 2'b10;	 rom[2][24][6] = 2'b10;	 rom[2][25][6] = 2'b10;	 rom[2][26][6] = 2'b10;	 rom[2][27][6] = 2'b01;	 rom[2][28][6] = 2'b01;	 rom[2][29][6] = 2'b10;	 rom[2][30][6] = 2'b10;	 rom[2][31][6] = 2'b00;	 rom[2][32][6] = 2'b00;	 rom[2][33][6] = 2'b00;	 rom[2][34][6] = 2'b00;	 rom[2][35][6] = 2'b00;	 rom[2][36][6] = 2'b00;	 rom[2][37][6] = 2'b00;	 rom[2][38][6] = 2'b00;	 rom[2][39][6] = 2'b00;
 rom[2][0][7] = 2'b10;	 rom[2][1][7] = 2'b10;	 rom[2][2][7] = 2'b10;	 rom[2][3][7] = 2'b10;	 rom[2][4][7] = 2'b10;	 rom[2][5][7] = 2'b10;	 rom[2][6][7] = 2'b10;	 rom[2][7][7] = 2'b10;	 rom[2][8][7] = 2'b10;	 rom[2][9][7] = 2'b10;	 rom[2][10][7] = 2'b10;	 rom[2][11][7] = 2'b10;	 rom[2][12][7] = 2'b10;	 rom[2][13][7] = 2'b10;	 rom[2][14][7] = 2'b10;	 rom[2][15][7] = 2'b10;	 rom[2][16][7] = 2'b10;	 rom[2][17][7] = 2'b10;	 rom[2][18][7] = 2'b10;	 rom[2][19][7] = 2'b10;	 rom[2][20][7] = 2'b10;	 rom[2][21][7] = 2'b10;	 rom[2][22][7] = 2'b10;	 rom[2][23][7] = 2'b10;	 rom[2][24][7] = 2'b10;	 rom[2][25][7] = 2'b10;	 rom[2][26][7] = 2'b10;	 rom[2][27][7] = 2'b10;	 rom[2][28][7] = 2'b01;	 rom[2][29][7] = 2'b10;	 rom[2][30][7] = 2'b10;	 rom[2][31][7] = 2'b00;	 rom[2][32][7] = 2'b00;	 rom[2][33][7] = 2'b00;	 rom[2][34][7] = 2'b00;	 rom[2][35][7] = 2'b00;	 rom[2][36][7] = 2'b00;	 rom[2][37][7] = 2'b00;	 rom[2][38][7] = 2'b00;	 rom[2][39][7] = 2'b00;
 rom[2][0][8] = 2'b10;	 rom[2][1][8] = 2'b11;	 rom[2][2][8] = 2'b11;	 rom[2][3][8] = 2'b11;	 rom[2][4][8] = 2'b11;	 rom[2][5][8] = 2'b11;	 rom[2][6][8] = 2'b11;	 rom[2][7][8] = 2'b11;	 rom[2][8][8] = 2'b11;	 rom[2][9][8] = 2'b11;	 rom[2][10][8] = 2'b11;	 rom[2][11][8] = 2'b11;	 rom[2][12][8] = 2'b11;	 rom[2][13][8] = 2'b11;	 rom[2][14][8] = 2'b11;	 rom[2][15][8] = 2'b11;	 rom[2][16][8] = 2'b10;	 rom[2][17][8] = 2'b10;	 rom[2][18][8] = 2'b10;	 rom[2][19][8] = 2'b10;	 rom[2][20][8] = 2'b01;	 rom[2][21][8] = 2'b01;	 rom[2][22][8] = 2'b10;	 rom[2][23][8] = 2'b01;	 rom[2][24][8] = 2'b01;	 rom[2][25][8] = 2'b10;	 rom[2][26][8] = 2'b10;	 rom[2][27][8] = 2'b10;	 rom[2][28][8] = 2'b10;	 rom[2][29][8] = 2'b10;	 rom[2][30][8] = 2'b10;	 rom[2][31][8] = 2'b10;	 rom[2][32][8] = 2'b10;	 rom[2][33][8] = 2'b10;	 rom[2][34][8] = 2'b00;	 rom[2][35][8] = 2'b00;	 rom[2][36][8] = 2'b00;	 rom[2][37][8] = 2'b00;	 rom[2][38][8] = 2'b00;	 rom[2][39][8] = 2'b00;
 rom[2][0][9] = 2'b10;	 rom[2][1][9] = 2'b11;	 rom[2][2][9] = 2'b11;	 rom[2][3][9] = 2'b11;	 rom[2][4][9] = 2'b11;	 rom[2][5][9] = 2'b11;	 rom[2][6][9] = 2'b11;	 rom[2][7][9] = 2'b11;	 rom[2][8][9] = 2'b11;	 rom[2][9][9] = 2'b11;	 rom[2][10][9] = 2'b11;	 rom[2][11][9] = 2'b11;	 rom[2][12][9] = 2'b11;	 rom[2][13][9] = 2'b11;	 rom[2][14][9] = 2'b11;	 rom[2][15][9] = 2'b10;	 rom[2][16][9] = 2'b10;	 rom[2][17][9] = 2'b01;	 rom[2][18][9] = 2'b01;	 rom[2][19][9] = 2'b01;	 rom[2][20][9] = 2'b01;	 rom[2][21][9] = 2'b01;	 rom[2][22][9] = 2'b01;	 rom[2][23][9] = 2'b01;	 rom[2][24][9] = 2'b01;	 rom[2][25][9] = 2'b01;	 rom[2][26][9] = 2'b01;	 rom[2][27][9] = 2'b10;	 rom[2][28][9] = 2'b10;	 rom[2][29][9] = 2'b10;	 rom[2][30][9] = 2'b10;	 rom[2][31][9] = 2'b10;	 rom[2][32][9] = 2'b10;	 rom[2][33][9] = 2'b10;	 rom[2][34][9] = 2'b10;	 rom[2][35][9] = 2'b10;	 rom[2][36][9] = 2'b00;	 rom[2][37][9] = 2'b00;	 rom[2][38][9] = 2'b00;	 rom[2][39][9] = 2'b00;
 rom[2][0][10] = 2'b10;	 rom[2][1][10] = 2'b10;	 rom[2][2][10] = 2'b10;	 rom[2][3][10] = 2'b10;	 rom[2][4][10] = 2'b10;	 rom[2][5][10] = 2'b10;	 rom[2][6][10] = 2'b10;	 rom[2][7][10] = 2'b10;	 rom[2][8][10] = 2'b10;	 rom[2][9][10] = 2'b10;	 rom[2][10][10] = 2'b10;	 rom[2][11][10] = 2'b10;	 rom[2][12][10] = 2'b10;	 rom[2][13][10] = 2'b10;	 rom[2][14][10] = 2'b10;	 rom[2][15][10] = 2'b10;	 rom[2][16][10] = 2'b01;	 rom[2][17][10] = 2'b01;	 rom[2][18][10] = 2'b01;	 rom[2][19][10] = 2'b01;	 rom[2][20][10] = 2'b01;	 rom[2][21][10] = 2'b01;	 rom[2][22][10] = 2'b01;	 rom[2][23][10] = 2'b01;	 rom[2][24][10] = 2'b01;	 rom[2][25][10] = 2'b01;	 rom[2][26][10] = 2'b01;	 rom[2][27][10] = 2'b01;	 rom[2][28][10] = 2'b10;	 rom[2][29][10] = 2'b10;	 rom[2][30][10] = 2'b10;	 rom[2][31][10] = 2'b10;	 rom[2][32][10] = 2'b10;	 rom[2][33][10] = 2'b10;	 rom[2][34][10] = 2'b10;	 rom[2][35][10] = 2'b10;	 rom[2][36][10] = 2'b10;	 rom[2][37][10] = 2'b10;	 rom[2][38][10] = 2'b00;	 rom[2][39][10] = 2'b00;
 rom[2][0][11] = 2'b10;	 rom[2][1][11] = 2'b10;	 rom[2][2][11] = 2'b00;	 rom[2][3][11] = 2'b00;	 rom[2][4][11] = 2'b00;	 rom[2][5][11] = 2'b00;	 rom[2][6][11] = 2'b00;	 rom[2][7][11] = 2'b00;	 rom[2][8][11] = 2'b00;	 rom[2][9][11] = 2'b00;	 rom[2][10][11] = 2'b00;	 rom[2][11][11] = 2'b00;	 rom[2][12][11] = 2'b00;	 rom[2][13][11] = 2'b10;	 rom[2][14][11] = 2'b10;	 rom[2][15][11] = 2'b01;	 rom[2][16][11] = 2'b01;	 rom[2][17][11] = 2'b01;	 rom[2][18][11] = 2'b01;	 rom[2][19][11] = 2'b01;	 rom[2][20][11] = 2'b01;	 rom[2][21][11] = 2'b01;	 rom[2][22][11] = 2'b01;	 rom[2][23][11] = 2'b01;	 rom[2][24][11] = 2'b01;	 rom[2][25][11] = 2'b01;	 rom[2][26][11] = 2'b01;	 rom[2][27][11] = 2'b01;	 rom[2][28][11] = 2'b01;	 rom[2][29][11] = 2'b10;	 rom[2][30][11] = 2'b10;	 rom[2][31][11] = 2'b10;	 rom[2][32][11] = 2'b10;	 rom[2][33][11] = 2'b10;	 rom[2][34][11] = 2'b11;	 rom[2][35][11] = 2'b11;	 rom[2][36][11] = 2'b11;	 rom[2][37][11] = 2'b10;	 rom[2][38][11] = 2'b00;	 rom[2][39][11] = 2'b00;
 rom[2][0][12] = 2'b00;	 rom[2][1][12] = 2'b00;	 rom[2][2][12] = 2'b00;	 rom[2][3][12] = 2'b00;	 rom[2][4][12] = 2'b00;	 rom[2][5][12] = 2'b00;	 rom[2][6][12] = 2'b00;	 rom[2][7][12] = 2'b00;	 rom[2][8][12] = 2'b00;	 rom[2][9][12] = 2'b00;	 rom[2][10][12] = 2'b00;	 rom[2][11][12] = 2'b10;	 rom[2][12][12] = 2'b10;	 rom[2][13][12] = 2'b10;	 rom[2][14][12] = 2'b01;	 rom[2][15][12] = 2'b01;	 rom[2][16][12] = 2'b01;	 rom[2][17][12] = 2'b01;	 rom[2][18][12] = 2'b01;	 rom[2][19][12] = 2'b01;	 rom[2][20][12] = 2'b01;	 rom[2][21][12] = 2'b01;	 rom[2][22][12] = 2'b01;	 rom[2][23][12] = 2'b01;	 rom[2][24][12] = 2'b01;	 rom[2][25][12] = 2'b01;	 rom[2][26][12] = 2'b01;	 rom[2][27][12] = 2'b01;	 rom[2][28][12] = 2'b01;	 rom[2][29][12] = 2'b01;	 rom[2][30][12] = 2'b10;	 rom[2][31][12] = 2'b10;	 rom[2][32][12] = 2'b10;	 rom[2][33][12] = 2'b11;	 rom[2][34][12] = 2'b11;	 rom[2][35][12] = 2'b11;	 rom[2][36][12] = 2'b11;	 rom[2][37][12] = 2'b10;	 rom[2][38][12] = 2'b00;	 rom[2][39][12] = 2'b00;
 rom[2][0][13] = 2'b00;	 rom[2][1][13] = 2'b00;	 rom[2][2][13] = 2'b00;	 rom[2][3][13] = 2'b00;	 rom[2][4][13] = 2'b00;	 rom[2][5][13] = 2'b00;	 rom[2][6][13] = 2'b00;	 rom[2][7][13] = 2'b00;	 rom[2][8][13] = 2'b10;	 rom[2][9][13] = 2'b10;	 rom[2][10][13] = 2'b10;	 rom[2][11][13] = 2'b10;	 rom[2][12][13] = 2'b10;	 rom[2][13][13] = 2'b01;	 rom[2][14][13] = 2'b01;	 rom[2][15][13] = 2'b01;	 rom[2][16][13] = 2'b01;	 rom[2][17][13] = 2'b01;	 rom[2][18][13] = 2'b01;	 rom[2][19][13] = 2'b01;	 rom[2][20][13] = 2'b01;	 rom[2][21][13] = 2'b01;	 rom[2][22][13] = 2'b01;	 rom[2][23][13] = 2'b01;	 rom[2][24][13] = 2'b01;	 rom[2][25][13] = 2'b01;	 rom[2][26][13] = 2'b01;	 rom[2][27][13] = 2'b01;	 rom[2][28][13] = 2'b01;	 rom[2][29][13] = 2'b01;	 rom[2][30][13] = 2'b10;	 rom[2][31][13] = 2'b11;	 rom[2][32][13] = 2'b11;	 rom[2][33][13] = 2'b11;	 rom[2][34][13] = 2'b11;	 rom[2][35][13] = 2'b11;	 rom[2][36][13] = 2'b11;	 rom[2][37][13] = 2'b10;	 rom[2][38][13] = 2'b00;	 rom[2][39][13] = 2'b00;
 rom[2][0][14] = 2'b00;	 rom[2][1][14] = 2'b00;	 rom[2][2][14] = 2'b00;	 rom[2][3][14] = 2'b00;	 rom[2][4][14] = 2'b00;	 rom[2][5][14] = 2'b00;	 rom[2][6][14] = 2'b00;	 rom[2][7][14] = 2'b10;	 rom[2][8][14] = 2'b10;	 rom[2][9][14] = 2'b11;	 rom[2][10][14] = 2'b10;	 rom[2][11][14] = 2'b10;	 rom[2][12][14] = 2'b01;	 rom[2][13][14] = 2'b01;	 rom[2][14][14] = 2'b01;	 rom[2][15][14] = 2'b01;	 rom[2][16][14] = 2'b01;	 rom[2][17][14] = 2'b01;	 rom[2][18][14] = 2'b01;	 rom[2][19][14] = 2'b01;	 rom[2][20][14] = 2'b01;	 rom[2][21][14] = 2'b01;	 rom[2][22][14] = 2'b01;	 rom[2][23][14] = 2'b01;	 rom[2][24][14] = 2'b01;	 rom[2][25][14] = 2'b01;	 rom[2][26][14] = 2'b01;	 rom[2][27][14] = 2'b01;	 rom[2][28][14] = 2'b01;	 rom[2][29][14] = 2'b01;	 rom[2][30][14] = 2'b10;	 rom[2][31][14] = 2'b11;	 rom[2][32][14] = 2'b11;	 rom[2][33][14] = 2'b11;	 rom[2][34][14] = 2'b11;	 rom[2][35][14] = 2'b11;	 rom[2][36][14] = 2'b11;	 rom[2][37][14] = 2'b10;	 rom[2][38][14] = 2'b00;	 rom[2][39][14] = 2'b00;
 rom[2][0][15] = 2'b00;	 rom[2][1][15] = 2'b00;	 rom[2][2][15] = 2'b00;	 rom[2][3][15] = 2'b00;	 rom[2][4][15] = 2'b00;	 rom[2][5][15] = 2'b00;	 rom[2][6][15] = 2'b10;	 rom[2][7][15] = 2'b10;	 rom[2][8][15] = 2'b11;	 rom[2][9][15] = 2'b11;	 rom[2][10][15] = 2'b10;	 rom[2][11][15] = 2'b10;	 rom[2][12][15] = 2'b01;	 rom[2][13][15] = 2'b01;	 rom[2][14][15] = 2'b01;	 rom[2][15][15] = 2'b01;	 rom[2][16][15] = 2'b01;	 rom[2][17][15] = 2'b01;	 rom[2][18][15] = 2'b01;	 rom[2][19][15] = 2'b01;	 rom[2][20][15] = 2'b01;	 rom[2][21][15] = 2'b01;	 rom[2][22][15] = 2'b01;	 rom[2][23][15] = 2'b01;	 rom[2][24][15] = 2'b01;	 rom[2][25][15] = 2'b01;	 rom[2][26][15] = 2'b01;	 rom[2][27][15] = 2'b01;	 rom[2][28][15] = 2'b01;	 rom[2][29][15] = 2'b01;	 rom[2][30][15] = 2'b10;	 rom[2][31][15] = 2'b10;	 rom[2][32][15] = 2'b10;	 rom[2][33][15] = 2'b10;	 rom[2][34][15] = 2'b11;	 rom[2][35][15] = 2'b11;	 rom[2][36][15] = 2'b11;	 rom[2][37][15] = 2'b10;	 rom[2][38][15] = 2'b00;	 rom[2][39][15] = 2'b00;
 rom[2][0][16] = 2'b00;	 rom[2][1][16] = 2'b00;	 rom[2][2][16] = 2'b00;	 rom[2][3][16] = 2'b00;	 rom[2][4][16] = 2'b00;	 rom[2][5][16] = 2'b00;	 rom[2][6][16] = 2'b10;	 rom[2][7][16] = 2'b11;	 rom[2][8][16] = 2'b11;	 rom[2][9][16] = 2'b11;	 rom[2][10][16] = 2'b10;	 rom[2][11][16] = 2'b10;	 rom[2][12][16] = 2'b01;	 rom[2][13][16] = 2'b01;	 rom[2][14][16] = 2'b01;	 rom[2][15][16] = 2'b01;	 rom[2][16][16] = 2'b01;	 rom[2][17][16] = 2'b01;	 rom[2][18][16] = 2'b01;	 rom[2][19][16] = 2'b01;	 rom[2][20][16] = 2'b01;	 rom[2][21][16] = 2'b01;	 rom[2][22][16] = 2'b01;	 rom[2][23][16] = 2'b01;	 rom[2][24][16] = 2'b01;	 rom[2][25][16] = 2'b01;	 rom[2][26][16] = 2'b01;	 rom[2][27][16] = 2'b01;	 rom[2][28][16] = 2'b01;	 rom[2][29][16] = 2'b01;	 rom[2][30][16] = 2'b01;	 rom[2][31][16] = 2'b10;	 rom[2][32][16] = 2'b10;	 rom[2][33][16] = 2'b10;	 rom[2][34][16] = 2'b11;	 rom[2][35][16] = 2'b11;	 rom[2][36][16] = 2'b11;	 rom[2][37][16] = 2'b10;	 rom[2][38][16] = 2'b00;	 rom[2][39][16] = 2'b00;
 rom[2][0][17] = 2'b00;	 rom[2][1][17] = 2'b00;	 rom[2][2][17] = 2'b00;	 rom[2][3][17] = 2'b00;	 rom[2][4][17] = 2'b00;	 rom[2][5][17] = 2'b00;	 rom[2][6][17] = 2'b10;	 rom[2][7][17] = 2'b11;	 rom[2][8][17] = 2'b11;	 rom[2][9][17] = 2'b11;	 rom[2][10][17] = 2'b10;	 rom[2][11][17] = 2'b10;	 rom[2][12][17] = 2'b01;	 rom[2][13][17] = 2'b01;	 rom[2][14][17] = 2'b01;	 rom[2][15][17] = 2'b01;	 rom[2][16][17] = 2'b01;	 rom[2][17][17] = 2'b01;	 rom[2][18][17] = 2'b01;	 rom[2][19][17] = 2'b01;	 rom[2][20][17] = 2'b01;	 rom[2][21][17] = 2'b01;	 rom[2][22][17] = 2'b01;	 rom[2][23][17] = 2'b01;	 rom[2][24][17] = 2'b01;	 rom[2][25][17] = 2'b01;	 rom[2][26][17] = 2'b01;	 rom[2][27][17] = 2'b01;	 rom[2][28][17] = 2'b01;	 rom[2][29][17] = 2'b01;	 rom[2][30][17] = 2'b01;	 rom[2][31][17] = 2'b10;	 rom[2][32][17] = 2'b10;	 rom[2][33][17] = 2'b10;	 rom[2][34][17] = 2'b11;	 rom[2][35][17] = 2'b10;	 rom[2][36][17] = 2'b11;	 rom[2][37][17] = 2'b10;	 rom[2][38][17] = 2'b00;	 rom[2][39][17] = 2'b00;
 rom[2][0][18] = 2'b00;	 rom[2][1][18] = 2'b00;	 rom[2][2][18] = 2'b00;	 rom[2][3][18] = 2'b00;	 rom[2][4][18] = 2'b00;	 rom[2][5][18] = 2'b00;	 rom[2][6][18] = 2'b10;	 rom[2][7][18] = 2'b11;	 rom[2][8][18] = 2'b11;	 rom[2][9][18] = 2'b11;	 rom[2][10][18] = 2'b10;	 rom[2][11][18] = 2'b10;	 rom[2][12][18] = 2'b01;	 rom[2][13][18] = 2'b01;	 rom[2][14][18] = 2'b01;	 rom[2][15][18] = 2'b01;	 rom[2][16][18] = 2'b01;	 rom[2][17][18] = 2'b01;	 rom[2][18][18] = 2'b01;	 rom[2][19][18] = 2'b01;	 rom[2][20][18] = 2'b01;	 rom[2][21][18] = 2'b01;	 rom[2][22][18] = 2'b01;	 rom[2][23][18] = 2'b01;	 rom[2][24][18] = 2'b01;	 rom[2][25][18] = 2'b01;	 rom[2][26][18] = 2'b01;	 rom[2][27][18] = 2'b01;	 rom[2][28][18] = 2'b01;	 rom[2][29][18] = 2'b01;	 rom[2][30][18] = 2'b01;	 rom[2][31][18] = 2'b10;	 rom[2][32][18] = 2'b10;	 rom[2][33][18] = 2'b10;	 rom[2][34][18] = 2'b11;	 rom[2][35][18] = 2'b10;	 rom[2][36][18] = 2'b11;	 rom[2][37][18] = 2'b10;	 rom[2][38][18] = 2'b00;	 rom[2][39][18] = 2'b00;
 rom[2][0][19] = 2'b00;	 rom[2][1][19] = 2'b00;	 rom[2][2][19] = 2'b00;	 rom[2][3][19] = 2'b00;	 rom[2][4][19] = 2'b00;	 rom[2][5][19] = 2'b00;	 rom[2][6][19] = 2'b10;	 rom[2][7][19] = 2'b11;	 rom[2][8][19] = 2'b11;	 rom[2][9][19] = 2'b11;	 rom[2][10][19] = 2'b10;	 rom[2][11][19] = 2'b10;	 rom[2][12][19] = 2'b01;	 rom[2][13][19] = 2'b01;	 rom[2][14][19] = 2'b01;	 rom[2][15][19] = 2'b01;	 rom[2][16][19] = 2'b01;	 rom[2][17][19] = 2'b01;	 rom[2][18][19] = 2'b01;	 rom[2][19][19] = 2'b01;	 rom[2][20][19] = 2'b01;	 rom[2][21][19] = 2'b01;	 rom[2][22][19] = 2'b01;	 rom[2][23][19] = 2'b01;	 rom[2][24][19] = 2'b01;	 rom[2][25][19] = 2'b01;	 rom[2][26][19] = 2'b01;	 rom[2][27][19] = 2'b01;	 rom[2][28][19] = 2'b01;	 rom[2][29][19] = 2'b01;	 rom[2][30][19] = 2'b01;	 rom[2][31][19] = 2'b10;	 rom[2][32][19] = 2'b10;	 rom[2][33][19] = 2'b10;	 rom[2][34][19] = 2'b11;	 rom[2][35][19] = 2'b10;	 rom[2][36][19] = 2'b11;	 rom[2][37][19] = 2'b10;	 rom[2][38][19] = 2'b00;	 rom[2][39][19] = 2'b00;
 rom[2][0][20] = 2'b00;	 rom[2][1][20] = 2'b00;	 rom[2][2][20] = 2'b00;	 rom[2][3][20] = 2'b00;	 rom[2][4][20] = 2'b00;	 rom[2][5][20] = 2'b00;	 rom[2][6][20] = 2'b10;	 rom[2][7][20] = 2'b10;	 rom[2][8][20] = 2'b11;	 rom[2][9][20] = 2'b11;	 rom[2][10][20] = 2'b10;	 rom[2][11][20] = 2'b10;	 rom[2][12][20] = 2'b01;	 rom[2][13][20] = 2'b01;	 rom[2][14][20] = 2'b01;	 rom[2][15][20] = 2'b01;	 rom[2][16][20] = 2'b01;	 rom[2][17][20] = 2'b01;	 rom[2][18][20] = 2'b01;	 rom[2][19][20] = 2'b01;	 rom[2][20][20] = 2'b01;	 rom[2][21][20] = 2'b01;	 rom[2][22][20] = 2'b01;	 rom[2][23][20] = 2'b01;	 rom[2][24][20] = 2'b01;	 rom[2][25][20] = 2'b01;	 rom[2][26][20] = 2'b01;	 rom[2][27][20] = 2'b01;	 rom[2][28][20] = 2'b01;	 rom[2][29][20] = 2'b01;	 rom[2][30][20] = 2'b01;	 rom[2][31][20] = 2'b10;	 rom[2][32][20] = 2'b10;	 rom[2][33][20] = 2'b10;	 rom[2][34][20] = 2'b11;	 rom[2][35][20] = 2'b10;	 rom[2][36][20] = 2'b11;	 rom[2][37][20] = 2'b10;	 rom[2][38][20] = 2'b00;	 rom[2][39][20] = 2'b00;
 rom[2][0][21] = 2'b00;	 rom[2][1][21] = 2'b00;	 rom[2][2][21] = 2'b00;	 rom[2][3][21] = 2'b00;	 rom[2][4][21] = 2'b00;	 rom[2][5][21] = 2'b00;	 rom[2][6][21] = 2'b00;	 rom[2][7][21] = 2'b10;	 rom[2][8][21] = 2'b10;	 rom[2][9][21] = 2'b10;	 rom[2][10][21] = 2'b10;	 rom[2][11][21] = 2'b10;	 rom[2][12][21] = 2'b01;	 rom[2][13][21] = 2'b01;	 rom[2][14][21] = 2'b01;	 rom[2][15][21] = 2'b01;	 rom[2][16][21] = 2'b01;	 rom[2][17][21] = 2'b01;	 rom[2][18][21] = 2'b01;	 rom[2][19][21] = 2'b01;	 rom[2][20][21] = 2'b01;	 rom[2][21][21] = 2'b01;	 rom[2][22][21] = 2'b01;	 rom[2][23][21] = 2'b01;	 rom[2][24][21] = 2'b01;	 rom[2][25][21] = 2'b01;	 rom[2][26][21] = 2'b01;	 rom[2][27][21] = 2'b01;	 rom[2][28][21] = 2'b01;	 rom[2][29][21] = 2'b01;	 rom[2][30][21] = 2'b01;	 rom[2][31][21] = 2'b10;	 rom[2][32][21] = 2'b10;	 rom[2][33][21] = 2'b10;	 rom[2][34][21] = 2'b11;	 rom[2][35][21] = 2'b10;	 rom[2][36][21] = 2'b11;	 rom[2][37][21] = 2'b10;	 rom[2][38][21] = 2'b00;	 rom[2][39][21] = 2'b00;
 rom[2][0][22] = 2'b00;	 rom[2][1][22] = 2'b00;	 rom[2][2][22] = 2'b00;	 rom[2][3][22] = 2'b00;	 rom[2][4][22] = 2'b00;	 rom[2][5][22] = 2'b00;	 rom[2][6][22] = 2'b00;	 rom[2][7][22] = 2'b00;	 rom[2][8][22] = 2'b00;	 rom[2][9][22] = 2'b00;	 rom[2][10][22] = 2'b10;	 rom[2][11][22] = 2'b10;	 rom[2][12][22] = 2'b01;	 rom[2][13][22] = 2'b01;	 rom[2][14][22] = 2'b01;	 rom[2][15][22] = 2'b01;	 rom[2][16][22] = 2'b01;	 rom[2][17][22] = 2'b01;	 rom[2][18][22] = 2'b01;	 rom[2][19][22] = 2'b01;	 rom[2][20][22] = 2'b01;	 rom[2][21][22] = 2'b01;	 rom[2][22][22] = 2'b01;	 rom[2][23][22] = 2'b01;	 rom[2][24][22] = 2'b01;	 rom[2][25][22] = 2'b01;	 rom[2][26][22] = 2'b01;	 rom[2][27][22] = 2'b01;	 rom[2][28][22] = 2'b01;	 rom[2][29][22] = 2'b01;	 rom[2][30][22] = 2'b01;	 rom[2][31][22] = 2'b10;	 rom[2][32][22] = 2'b10;	 rom[2][33][22] = 2'b10;	 rom[2][34][22] = 2'b11;	 rom[2][35][22] = 2'b10;	 rom[2][36][22] = 2'b11;	 rom[2][37][22] = 2'b10;	 rom[2][38][22] = 2'b00;	 rom[2][39][22] = 2'b00;
 rom[2][0][23] = 2'b00;	 rom[2][1][23] = 2'b00;	 rom[2][2][23] = 2'b00;	 rom[2][3][23] = 2'b00;	 rom[2][4][23] = 2'b00;	 rom[2][5][23] = 2'b00;	 rom[2][6][23] = 2'b00;	 rom[2][7][23] = 2'b00;	 rom[2][8][23] = 2'b00;	 rom[2][9][23] = 2'b10;	 rom[2][10][23] = 2'b10;	 rom[2][11][23] = 2'b10;	 rom[2][12][23] = 2'b01;	 rom[2][13][23] = 2'b01;	 rom[2][14][23] = 2'b01;	 rom[2][15][23] = 2'b01;	 rom[2][16][23] = 2'b01;	 rom[2][17][23] = 2'b01;	 rom[2][18][23] = 2'b01;	 rom[2][19][23] = 2'b01;	 rom[2][20][23] = 2'b01;	 rom[2][21][23] = 2'b01;	 rom[2][22][23] = 2'b01;	 rom[2][23][23] = 2'b01;	 rom[2][24][23] = 2'b01;	 rom[2][25][23] = 2'b01;	 rom[2][26][23] = 2'b01;	 rom[2][27][23] = 2'b01;	 rom[2][28][23] = 2'b01;	 rom[2][29][23] = 2'b01;	 rom[2][30][23] = 2'b01;	 rom[2][31][23] = 2'b10;	 rom[2][32][23] = 2'b10;	 rom[2][33][23] = 2'b10;	 rom[2][34][23] = 2'b11;	 rom[2][35][23] = 2'b11;	 rom[2][36][23] = 2'b11;	 rom[2][37][23] = 2'b10;	 rom[2][38][23] = 2'b00;	 rom[2][39][23] = 2'b00;
 rom[2][0][24] = 2'b00;	 rom[2][1][24] = 2'b00;	 rom[2][2][24] = 2'b00;	 rom[2][3][24] = 2'b00;	 rom[2][4][24] = 2'b00;	 rom[2][5][24] = 2'b00;	 rom[2][6][24] = 2'b00;	 rom[2][7][24] = 2'b00;	 rom[2][8][24] = 2'b10;	 rom[2][9][24] = 2'b10;	 rom[2][10][24] = 2'b10;	 rom[2][11][24] = 2'b10;	 rom[2][12][24] = 2'b01;	 rom[2][13][24] = 2'b01;	 rom[2][14][24] = 2'b01;	 rom[2][15][24] = 2'b01;	 rom[2][16][24] = 2'b01;	 rom[2][17][24] = 2'b01;	 rom[2][18][24] = 2'b01;	 rom[2][19][24] = 2'b01;	 rom[2][20][24] = 2'b01;	 rom[2][21][24] = 2'b01;	 rom[2][22][24] = 2'b01;	 rom[2][23][24] = 2'b01;	 rom[2][24][24] = 2'b01;	 rom[2][25][24] = 2'b01;	 rom[2][26][24] = 2'b01;	 rom[2][27][24] = 2'b01;	 rom[2][28][24] = 2'b01;	 rom[2][29][24] = 2'b01;	 rom[2][30][24] = 2'b10;	 rom[2][31][24] = 2'b10;	 rom[2][32][24] = 2'b10;	 rom[2][33][24] = 2'b10;	 rom[2][34][24] = 2'b11;	 rom[2][35][24] = 2'b11;	 rom[2][36][24] = 2'b11;	 rom[2][37][24] = 2'b10;	 rom[2][38][24] = 2'b00;	 rom[2][39][24] = 2'b00;
 rom[2][0][25] = 2'b00;	 rom[2][1][25] = 2'b00;	 rom[2][2][25] = 2'b00;	 rom[2][3][25] = 2'b00;	 rom[2][4][25] = 2'b00;	 rom[2][5][25] = 2'b00;	 rom[2][6][25] = 2'b00;	 rom[2][7][25] = 2'b10;	 rom[2][8][25] = 2'b10;	 rom[2][9][25] = 2'b11;	 rom[2][10][25] = 2'b10;	 rom[2][11][25] = 2'b10;	 rom[2][12][25] = 2'b01;	 rom[2][13][25] = 2'b01;	 rom[2][14][25] = 2'b01;	 rom[2][15][25] = 2'b01;	 rom[2][16][25] = 2'b01;	 rom[2][17][25] = 2'b01;	 rom[2][18][25] = 2'b01;	 rom[2][19][25] = 2'b01;	 rom[2][20][25] = 2'b01;	 rom[2][21][25] = 2'b01;	 rom[2][22][25] = 2'b01;	 rom[2][23][25] = 2'b01;	 rom[2][24][25] = 2'b01;	 rom[2][25][25] = 2'b01;	 rom[2][26][25] = 2'b01;	 rom[2][27][25] = 2'b01;	 rom[2][28][25] = 2'b01;	 rom[2][29][25] = 2'b01;	 rom[2][30][25] = 2'b10;	 rom[2][31][25] = 2'b11;	 rom[2][32][25] = 2'b11;	 rom[2][33][25] = 2'b11;	 rom[2][34][25] = 2'b11;	 rom[2][35][25] = 2'b11;	 rom[2][36][25] = 2'b11;	 rom[2][37][25] = 2'b10;	 rom[2][38][25] = 2'b00;	 rom[2][39][25] = 2'b00;
 rom[2][0][26] = 2'b00;	 rom[2][1][26] = 2'b00;	 rom[2][2][26] = 2'b00;	 rom[2][3][26] = 2'b00;	 rom[2][4][26] = 2'b00;	 rom[2][5][26] = 2'b00;	 rom[2][6][26] = 2'b00;	 rom[2][7][26] = 2'b10;	 rom[2][8][26] = 2'b11;	 rom[2][9][26] = 2'b11;	 rom[2][10][26] = 2'b11;	 rom[2][11][26] = 2'b10;	 rom[2][12][26] = 2'b10;	 rom[2][13][26] = 2'b01;	 rom[2][14][26] = 2'b01;	 rom[2][15][26] = 2'b01;	 rom[2][16][26] = 2'b01;	 rom[2][17][26] = 2'b01;	 rom[2][18][26] = 2'b01;	 rom[2][19][26] = 2'b01;	 rom[2][20][26] = 2'b01;	 rom[2][21][26] = 2'b01;	 rom[2][22][26] = 2'b01;	 rom[2][23][26] = 2'b01;	 rom[2][24][26] = 2'b01;	 rom[2][25][26] = 2'b01;	 rom[2][26][26] = 2'b01;	 rom[2][27][26] = 2'b01;	 rom[2][28][26] = 2'b01;	 rom[2][29][26] = 2'b01;	 rom[2][30][26] = 2'b10;	 rom[2][31][26] = 2'b11;	 rom[2][32][26] = 2'b11;	 rom[2][33][26] = 2'b11;	 rom[2][34][26] = 2'b11;	 rom[2][35][26] = 2'b11;	 rom[2][36][26] = 2'b11;	 rom[2][37][26] = 2'b10;	 rom[2][38][26] = 2'b00;	 rom[2][39][26] = 2'b00;
 rom[2][0][27] = 2'b00;	 rom[2][1][27] = 2'b00;	 rom[2][2][27] = 2'b00;	 rom[2][3][27] = 2'b00;	 rom[2][4][27] = 2'b00;	 rom[2][5][27] = 2'b00;	 rom[2][6][27] = 2'b00;	 rom[2][7][27] = 2'b10;	 rom[2][8][27] = 2'b11;	 rom[2][9][27] = 2'b11;	 rom[2][10][27] = 2'b11;	 rom[2][11][27] = 2'b10;	 rom[2][12][27] = 2'b10;	 rom[2][13][27] = 2'b10;	 rom[2][14][27] = 2'b01;	 rom[2][15][27] = 2'b01;	 rom[2][16][27] = 2'b01;	 rom[2][17][27] = 2'b01;	 rom[2][18][27] = 2'b01;	 rom[2][19][27] = 2'b01;	 rom[2][20][27] = 2'b01;	 rom[2][21][27] = 2'b01;	 rom[2][22][27] = 2'b01;	 rom[2][23][27] = 2'b01;	 rom[2][24][27] = 2'b01;	 rom[2][25][27] = 2'b01;	 rom[2][26][27] = 2'b01;	 rom[2][27][27] = 2'b01;	 rom[2][28][27] = 2'b01;	 rom[2][29][27] = 2'b01;	 rom[2][30][27] = 2'b10;	 rom[2][31][27] = 2'b10;	 rom[2][32][27] = 2'b10;	 rom[2][33][27] = 2'b11;	 rom[2][34][27] = 2'b11;	 rom[2][35][27] = 2'b11;	 rom[2][36][27] = 2'b11;	 rom[2][37][27] = 2'b10;	 rom[2][38][27] = 2'b00;	 rom[2][39][27] = 2'b00;
 rom[2][0][28] = 2'b00;	 rom[2][1][28] = 2'b00;	 rom[2][2][28] = 2'b00;	 rom[2][3][28] = 2'b00;	 rom[2][4][28] = 2'b00;	 rom[2][5][28] = 2'b00;	 rom[2][6][28] = 2'b00;	 rom[2][7][28] = 2'b10;	 rom[2][8][28] = 2'b11;	 rom[2][9][28] = 2'b11;	 rom[2][10][28] = 2'b11;	 rom[2][11][28] = 2'b11;	 rom[2][12][28] = 2'b11;	 rom[2][13][28] = 2'b10;	 rom[2][14][28] = 2'b10;	 rom[2][15][28] = 2'b01;	 rom[2][16][28] = 2'b01;	 rom[2][17][28] = 2'b01;	 rom[2][18][28] = 2'b01;	 rom[2][19][28] = 2'b01;	 rom[2][20][28] = 2'b01;	 rom[2][21][28] = 2'b01;	 rom[2][22][28] = 2'b01;	 rom[2][23][28] = 2'b01;	 rom[2][24][28] = 2'b01;	 rom[2][25][28] = 2'b01;	 rom[2][26][28] = 2'b01;	 rom[2][27][28] = 2'b01;	 rom[2][28][28] = 2'b01;	 rom[2][29][28] = 2'b10;	 rom[2][30][28] = 2'b10;	 rom[2][31][28] = 2'b10;	 rom[2][32][28] = 2'b10;	 rom[2][33][28] = 2'b10;	 rom[2][34][28] = 2'b11;	 rom[2][35][28] = 2'b11;	 rom[2][36][28] = 2'b11;	 rom[2][37][28] = 2'b10;	 rom[2][38][28] = 2'b00;	 rom[2][39][28] = 2'b00;
 rom[2][0][29] = 2'b00;	 rom[2][1][29] = 2'b00;	 rom[2][2][29] = 2'b00;	 rom[2][3][29] = 2'b00;	 rom[2][4][29] = 2'b00;	 rom[2][5][29] = 2'b00;	 rom[2][6][29] = 2'b00;	 rom[2][7][29] = 2'b10;	 rom[2][8][29] = 2'b11;	 rom[2][9][29] = 2'b11;	 rom[2][10][29] = 2'b11;	 rom[2][11][29] = 2'b11;	 rom[2][12][29] = 2'b11;	 rom[2][13][29] = 2'b10;	 rom[2][14][29] = 2'b10;	 rom[2][15][29] = 2'b10;	 rom[2][16][29] = 2'b01;	 rom[2][17][29] = 2'b01;	 rom[2][18][29] = 2'b01;	 rom[2][19][29] = 2'b01;	 rom[2][20][29] = 2'b01;	 rom[2][21][29] = 2'b01;	 rom[2][22][29] = 2'b01;	 rom[2][23][29] = 2'b01;	 rom[2][24][29] = 2'b01;	 rom[2][25][29] = 2'b01;	 rom[2][26][29] = 2'b01;	 rom[2][27][29] = 2'b01;	 rom[2][28][29] = 2'b10;	 rom[2][29][29] = 2'b10;	 rom[2][30][29] = 2'b10;	 rom[2][31][29] = 2'b10;	 rom[2][32][29] = 2'b10;	 rom[2][33][29] = 2'b10;	 rom[2][34][29] = 2'b10;	 rom[2][35][29] = 2'b10;	 rom[2][36][29] = 2'b10;	 rom[2][37][29] = 2'b10;	 rom[2][38][29] = 2'b00;	 rom[2][39][29] = 2'b00;
 rom[2][0][30] = 2'b00;	 rom[2][1][30] = 2'b00;	 rom[2][2][30] = 2'b00;	 rom[2][3][30] = 2'b00;	 rom[2][4][30] = 2'b00;	 rom[2][5][30] = 2'b00;	 rom[2][6][30] = 2'b00;	 rom[2][7][30] = 2'b10;	 rom[2][8][30] = 2'b10;	 rom[2][9][30] = 2'b11;	 rom[2][10][30] = 2'b11;	 rom[2][11][30] = 2'b11;	 rom[2][12][30] = 2'b11;	 rom[2][13][30] = 2'b11;	 rom[2][14][30] = 2'b10;	 rom[2][15][30] = 2'b10;	 rom[2][16][30] = 2'b10;	 rom[2][17][30] = 2'b01;	 rom[2][18][30] = 2'b01;	 rom[2][19][30] = 2'b01;	 rom[2][20][30] = 2'b01;	 rom[2][21][30] = 2'b01;	 rom[2][22][30] = 2'b01;	 rom[2][23][30] = 2'b01;	 rom[2][24][30] = 2'b01;	 rom[2][25][30] = 2'b01;	 rom[2][26][30] = 2'b01;	 rom[2][27][30] = 2'b10;	 rom[2][28][30] = 2'b10;	 rom[2][29][30] = 2'b10;	 rom[2][30][30] = 2'b10;	 rom[2][31][30] = 2'b10;	 rom[2][32][30] = 2'b10;	 rom[2][33][30] = 2'b10;	 rom[2][34][30] = 2'b10;	 rom[2][35][30] = 2'b10;	 rom[2][36][30] = 2'b00;	 rom[2][37][30] = 2'b00;	 rom[2][38][30] = 2'b00;	 rom[2][39][30] = 2'b00;
 rom[2][0][31] = 2'b00;	 rom[2][1][31] = 2'b00;	 rom[2][2][31] = 2'b00;	 rom[2][3][31] = 2'b00;	 rom[2][4][31] = 2'b00;	 rom[2][5][31] = 2'b00;	 rom[2][6][31] = 2'b00;	 rom[2][7][31] = 2'b00;	 rom[2][8][31] = 2'b10;	 rom[2][9][31] = 2'b10;	 rom[2][10][31] = 2'b11;	 rom[2][11][31] = 2'b11;	 rom[2][12][31] = 2'b11;	 rom[2][13][31] = 2'b11;	 rom[2][14][31] = 2'b11;	 rom[2][15][31] = 2'b10;	 rom[2][16][31] = 2'b10;	 rom[2][17][31] = 2'b10;	 rom[2][18][31] = 2'b10;	 rom[2][19][31] = 2'b10;	 rom[2][20][31] = 2'b01;	 rom[2][21][31] = 2'b01;	 rom[2][22][31] = 2'b01;	 rom[2][23][31] = 2'b01;	 rom[2][24][31] = 2'b01;	 rom[2][25][31] = 2'b01;	 rom[2][26][31] = 2'b10;	 rom[2][27][31] = 2'b10;	 rom[2][28][31] = 2'b10;	 rom[2][29][31] = 2'b10;	 rom[2][30][31] = 2'b10;	 rom[2][31][31] = 2'b10;	 rom[2][32][31] = 2'b10;	 rom[2][33][31] = 2'b10;	 rom[2][34][31] = 2'b00;	 rom[2][35][31] = 2'b00;	 rom[2][36][31] = 2'b00;	 rom[2][37][31] = 2'b00;	 rom[2][38][31] = 2'b00;	 rom[2][39][31] = 2'b00;
 rom[2][0][32] = 2'b00;	 rom[2][1][32] = 2'b00;	 rom[2][2][32] = 2'b00;	 rom[2][3][32] = 2'b00;	 rom[2][4][32] = 2'b00;	 rom[2][5][32] = 2'b00;	 rom[2][6][32] = 2'b00;	 rom[2][7][32] = 2'b00;	 rom[2][8][32] = 2'b00;	 rom[2][9][32] = 2'b10;	 rom[2][10][32] = 2'b10;	 rom[2][11][32] = 2'b10;	 rom[2][12][32] = 2'b10;	 rom[2][13][32] = 2'b10;	 rom[2][14][32] = 2'b10;	 rom[2][15][32] = 2'b10;	 rom[2][16][32] = 2'b00;	 rom[2][17][32] = 2'b10;	 rom[2][18][32] = 2'b10;	 rom[2][19][32] = 2'b10;	 rom[2][20][32] = 2'b10;	 rom[2][21][32] = 2'b10;	 rom[2][22][32] = 2'b10;	 rom[2][23][32] = 2'b10;	 rom[2][24][32] = 2'b10;	 rom[2][25][32] = 2'b10;	 rom[2][26][32] = 2'b10;	 rom[2][27][32] = 2'b10;	 rom[2][28][32] = 2'b01;	 rom[2][29][32] = 2'b10;	 rom[2][30][32] = 2'b10;	 rom[2][31][32] = 2'b00;	 rom[2][32][32] = 2'b00;	 rom[2][33][32] = 2'b00;	 rom[2][34][32] = 2'b00;	 rom[2][35][32] = 2'b00;	 rom[2][36][32] = 2'b00;	 rom[2][37][32] = 2'b00;	 rom[2][38][32] = 2'b00;	 rom[2][39][32] = 2'b00;
 rom[2][0][33] = 2'b00;	 rom[2][1][33] = 2'b00;	 rom[2][2][33] = 2'b00;	 rom[2][3][33] = 2'b00;	 rom[2][4][33] = 2'b00;	 rom[2][5][33] = 2'b00;	 rom[2][6][33] = 2'b00;	 rom[2][7][33] = 2'b00;	 rom[2][8][33] = 2'b00;	 rom[2][9][33] = 2'b00;	 rom[2][10][33] = 2'b00;	 rom[2][11][33] = 2'b00;	 rom[2][12][33] = 2'b00;	 rom[2][13][33] = 2'b00;	 rom[2][14][33] = 2'b00;	 rom[2][15][33] = 2'b00;	 rom[2][16][33] = 2'b00;	 rom[2][17][33] = 2'b10;	 rom[2][18][33] = 2'b10;	 rom[2][19][33] = 2'b10;	 rom[2][20][33] = 2'b10;	 rom[2][21][33] = 2'b10;	 rom[2][22][33] = 2'b10;	 rom[2][23][33] = 2'b10;	 rom[2][24][33] = 2'b10;	 rom[2][25][33] = 2'b10;	 rom[2][26][33] = 2'b10;	 rom[2][27][33] = 2'b01;	 rom[2][28][33] = 2'b01;	 rom[2][29][33] = 2'b10;	 rom[2][30][33] = 2'b10;	 rom[2][31][33] = 2'b00;	 rom[2][32][33] = 2'b00;	 rom[2][33][33] = 2'b00;	 rom[2][34][33] = 2'b00;	 rom[2][35][33] = 2'b00;	 rom[2][36][33] = 2'b00;	 rom[2][37][33] = 2'b00;	 rom[2][38][33] = 2'b00;	 rom[2][39][33] = 2'b00;
 rom[2][0][34] = 2'b00;	 rom[2][1][34] = 2'b00;	 rom[2][2][34] = 2'b00;	 rom[2][3][34] = 2'b00;	 rom[2][4][34] = 2'b00;	 rom[2][5][34] = 2'b00;	 rom[2][6][34] = 2'b00;	 rom[2][7][34] = 2'b00;	 rom[2][8][34] = 2'b00;	 rom[2][9][34] = 2'b00;	 rom[2][10][34] = 2'b00;	 rom[2][11][34] = 2'b00;	 rom[2][12][34] = 2'b00;	 rom[2][13][34] = 2'b00;	 rom[2][14][34] = 2'b00;	 rom[2][15][34] = 2'b00;	 rom[2][16][34] = 2'b00;	 rom[2][17][34] = 2'b00;	 rom[2][18][34] = 2'b10;	 rom[2][19][34] = 2'b01;	 rom[2][20][34] = 2'b01;	 rom[2][21][34] = 2'b01;	 rom[2][22][34] = 2'b01;	 rom[2][23][34] = 2'b01;	 rom[2][24][34] = 2'b01;	 rom[2][25][34] = 2'b01;	 rom[2][26][34] = 2'b01;	 rom[2][27][34] = 2'b01;	 rom[2][28][34] = 2'b01;	 rom[2][29][34] = 2'b10;	 rom[2][30][34] = 2'b10;	 rom[2][31][34] = 2'b00;	 rom[2][32][34] = 2'b00;	 rom[2][33][34] = 2'b00;	 rom[2][34][34] = 2'b00;	 rom[2][35][34] = 2'b00;	 rom[2][36][34] = 2'b00;	 rom[2][37][34] = 2'b00;	 rom[2][38][34] = 2'b00;	 rom[2][39][34] = 2'b00;
 rom[2][0][35] = 2'b00;	 rom[2][1][35] = 2'b00;	 rom[2][2][35] = 2'b00;	 rom[2][3][35] = 2'b00;	 rom[2][4][35] = 2'b00;	 rom[2][5][35] = 2'b00;	 rom[2][6][35] = 2'b00;	 rom[2][7][35] = 2'b00;	 rom[2][8][35] = 2'b00;	 rom[2][9][35] = 2'b00;	 rom[2][10][35] = 2'b00;	 rom[2][11][35] = 2'b00;	 rom[2][12][35] = 2'b00;	 rom[2][13][35] = 2'b00;	 rom[2][14][35] = 2'b00;	 rom[2][15][35] = 2'b00;	 rom[2][16][35] = 2'b00;	 rom[2][17][35] = 2'b00;	 rom[2][18][35] = 2'b10;	 rom[2][19][35] = 2'b10;	 rom[2][20][35] = 2'b01;	 rom[2][21][35] = 2'b01;	 rom[2][22][35] = 2'b01;	 rom[2][23][35] = 2'b01;	 rom[2][24][35] = 2'b01;	 rom[2][25][35] = 2'b01;	 rom[2][26][35] = 2'b01;	 rom[2][27][35] = 2'b01;	 rom[2][28][35] = 2'b01;	 rom[2][29][35] = 2'b10;	 rom[2][30][35] = 2'b10;	 rom[2][31][35] = 2'b00;	 rom[2][32][35] = 2'b00;	 rom[2][33][35] = 2'b00;	 rom[2][34][35] = 2'b00;	 rom[2][35][35] = 2'b00;	 rom[2][36][35] = 2'b00;	 rom[2][37][35] = 2'b00;	 rom[2][38][35] = 2'b00;	 rom[2][39][35] = 2'b00;
 rom[2][0][36] = 2'b00;	 rom[2][1][36] = 2'b00;	 rom[2][2][36] = 2'b00;	 rom[2][3][36] = 2'b00;	 rom[2][4][36] = 2'b00;	 rom[2][5][36] = 2'b00;	 rom[2][6][36] = 2'b00;	 rom[2][7][36] = 2'b00;	 rom[2][8][36] = 2'b00;	 rom[2][9][36] = 2'b00;	 rom[2][10][36] = 2'b00;	 rom[2][11][36] = 2'b00;	 rom[2][12][36] = 2'b00;	 rom[2][13][36] = 2'b00;	 rom[2][14][36] = 2'b00;	 rom[2][15][36] = 2'b00;	 rom[2][16][36] = 2'b00;	 rom[2][17][36] = 2'b00;	 rom[2][18][36] = 2'b00;	 rom[2][19][36] = 2'b10;	 rom[2][20][36] = 2'b10;	 rom[2][21][36] = 2'b01;	 rom[2][22][36] = 2'b01;	 rom[2][23][36] = 2'b01;	 rom[2][24][36] = 2'b01;	 rom[2][25][36] = 2'b01;	 rom[2][26][36] = 2'b01;	 rom[2][27][36] = 2'b01;	 rom[2][28][36] = 2'b10;	 rom[2][29][36] = 2'b10;	 rom[2][30][36] = 2'b00;	 rom[2][31][36] = 2'b00;	 rom[2][32][36] = 2'b00;	 rom[2][33][36] = 2'b00;	 rom[2][34][36] = 2'b00;	 rom[2][35][36] = 2'b00;	 rom[2][36][36] = 2'b00;	 rom[2][37][36] = 2'b00;	 rom[2][38][36] = 2'b00;	 rom[2][39][36] = 2'b00;
 rom[2][0][37] = 2'b00;	 rom[2][1][37] = 2'b00;	 rom[2][2][37] = 2'b00;	 rom[2][3][37] = 2'b00;	 rom[2][4][37] = 2'b00;	 rom[2][5][37] = 2'b00;	 rom[2][6][37] = 2'b00;	 rom[2][7][37] = 2'b00;	 rom[2][8][37] = 2'b00;	 rom[2][9][37] = 2'b00;	 rom[2][10][37] = 2'b00;	 rom[2][11][37] = 2'b00;	 rom[2][12][37] = 2'b00;	 rom[2][13][37] = 2'b00;	 rom[2][14][37] = 2'b00;	 rom[2][15][37] = 2'b00;	 rom[2][16][37] = 2'b00;	 rom[2][17][37] = 2'b00;	 rom[2][18][37] = 2'b00;	 rom[2][19][37] = 2'b10;	 rom[2][20][37] = 2'b10;	 rom[2][21][37] = 2'b10;	 rom[2][22][37] = 2'b10;	 rom[2][23][37] = 2'b10;	 rom[2][24][37] = 2'b10;	 rom[2][25][37] = 2'b10;	 rom[2][26][37] = 2'b10;	 rom[2][27][37] = 2'b10;	 rom[2][28][37] = 2'b10;	 rom[2][29][37] = 2'b00;	 rom[2][30][37] = 2'b00;	 rom[2][31][37] = 2'b00;	 rom[2][32][37] = 2'b00;	 rom[2][33][37] = 2'b00;	 rom[2][34][37] = 2'b00;	 rom[2][35][37] = 2'b00;	 rom[2][36][37] = 2'b00;	 rom[2][37][37] = 2'b00;	 rom[2][38][37] = 2'b00;	 rom[2][39][37] = 2'b00;
 rom[2][0][38] = 2'b00;	 rom[2][1][38] = 2'b00;	 rom[2][2][38] = 2'b00;	 rom[2][3][38] = 2'b00;	 rom[2][4][38] = 2'b00;	 rom[2][5][38] = 2'b00;	 rom[2][6][38] = 2'b00;	 rom[2][7][38] = 2'b00;	 rom[2][8][38] = 2'b00;	 rom[2][9][38] = 2'b00;	 rom[2][10][38] = 2'b00;	 rom[2][11][38] = 2'b00;	 rom[2][12][38] = 2'b00;	 rom[2][13][38] = 2'b00;	 rom[2][14][38] = 2'b00;	 rom[2][15][38] = 2'b00;	 rom[2][16][38] = 2'b00;	 rom[2][17][38] = 2'b00;	 rom[2][18][38] = 2'b00;	 rom[2][19][38] = 2'b00;	 rom[2][20][38] = 2'b00;	 rom[2][21][38] = 2'b00;	 rom[2][22][38] = 2'b00;	 rom[2][23][38] = 2'b00;	 rom[2][24][38] = 2'b00;	 rom[2][25][38] = 2'b00;	 rom[2][26][38] = 2'b00;	 rom[2][27][38] = 2'b00;	 rom[2][28][38] = 2'b00;	 rom[2][29][38] = 2'b00;	 rom[2][30][38] = 2'b00;	 rom[2][31][38] = 2'b00;	 rom[2][32][38] = 2'b00;	 rom[2][33][38] = 2'b00;	 rom[2][34][38] = 2'b00;	 rom[2][35][38] = 2'b00;	 rom[2][36][38] = 2'b00;	 rom[2][37][38] = 2'b00;	 rom[2][38][38] = 2'b00;	 rom[2][39][38] = 2'b00;
 rom[2][0][39] = 2'b00;	 rom[2][1][39] = 2'b00;	 rom[2][2][39] = 2'b00;	 rom[2][3][39] = 2'b00;	 rom[2][4][39] = 2'b00;	 rom[2][5][39] = 2'b00;	 rom[2][6][39] = 2'b00;	 rom[2][7][39] = 2'b00;	 rom[2][8][39] = 2'b00;	 rom[2][9][39] = 2'b00;	 rom[2][10][39] = 2'b00;	 rom[2][11][39] = 2'b00;	 rom[2][12][39] = 2'b00;	 rom[2][13][39] = 2'b00;	 rom[2][14][39] = 2'b00;	 rom[2][15][39] = 2'b00;	 rom[2][16][39] = 2'b00;	 rom[2][17][39] = 2'b00;	 rom[2][18][39] = 2'b00;	 rom[2][19][39] = 2'b00;	 rom[2][20][39] = 2'b00;	 rom[2][21][39] = 2'b00;	 rom[2][22][39] = 2'b00;	 rom[2][23][39] = 2'b00;	 rom[2][24][39] = 2'b00;	 rom[2][25][39] = 2'b00;	 rom[2][26][39] = 2'b00;	 rom[2][27][39] = 2'b00;	 rom[2][28][39] = 2'b00;	 rom[2][29][39] = 2'b00;	 rom[2][30][39] = 2'b00;	 rom[2][31][39] = 2'b00;	 rom[2][32][39] = 2'b00;	 rom[2][33][39] = 2'b00;	 rom[2][34][39] = 2'b00;	 rom[2][35][39] = 2'b00;	 rom[2][36][39] = 2'b00;	 rom[2][37][39] = 2'b00;	 rom[2][38][39] = 2'b00;	 rom[2][39][39] = 2'b00;

//right

 rom[3][0][0] = 2'b00;	 rom[3][1][0] = 2'b00;	 rom[3][2][0] = 2'b00;	 rom[3][3][0] = 2'b00;	 rom[3][4][0] = 2'b00;	 rom[3][5][0] = 2'b00;	 rom[3][6][0] = 2'b00;	 rom[3][7][0] = 2'b00;	 rom[3][8][0] = 2'b00;	 rom[3][9][0] = 2'b00;	 rom[3][10][0] = 2'b00;	 rom[3][11][0] = 2'b00;	 rom[3][12][0] = 2'b00;	 rom[3][13][0] = 2'b00;	 rom[3][14][0] = 2'b00;	 rom[3][15][0] = 2'b00;	 rom[3][16][0] = 2'b00;	 rom[3][17][0] = 2'b00;	 rom[3][18][0] = 2'b00;	 rom[3][19][0] = 2'b00;	 rom[3][20][0] = 2'b00;	 rom[3][21][0] = 2'b00;	 rom[3][22][0] = 2'b00;	 rom[3][23][0] = 2'b00;	 rom[3][24][0] = 2'b00;	 rom[3][25][0] = 2'b00;	 rom[3][26][0] = 2'b00;	 rom[3][27][0] = 2'b00;	 rom[3][28][0] = 2'b00;	 rom[3][29][0] = 2'b00;	 rom[3][30][0] = 2'b00;	 rom[3][31][0] = 2'b00;	 rom[3][32][0] = 2'b00;	 rom[3][33][0] = 2'b00;	 rom[3][34][0] = 2'b00;	 rom[3][35][0] = 2'b00;	 rom[3][36][0] = 2'b00;	 rom[3][37][0] = 2'b00;	 rom[3][38][0] = 2'b00;	 rom[3][39][0] = 2'b00;
 rom[3][0][1] = 2'b00;	 rom[3][1][1] = 2'b00;	 rom[3][2][1] = 2'b00;	 rom[3][3][1] = 2'b00;	 rom[3][4][1] = 2'b00;	 rom[3][5][1] = 2'b00;	 rom[3][6][1] = 2'b00;	 rom[3][7][1] = 2'b00;	 rom[3][8][1] = 2'b00;	 rom[3][9][1] = 2'b00;	 rom[3][10][1] = 2'b00;	 rom[3][11][1] = 2'b00;	 rom[3][12][1] = 2'b00;	 rom[3][13][1] = 2'b00;	 rom[3][14][1] = 2'b00;	 rom[3][15][1] = 2'b00;	 rom[3][16][1] = 2'b00;	 rom[3][17][1] = 2'b00;	 rom[3][18][1] = 2'b00;	 rom[3][19][1] = 2'b00;	 rom[3][20][1] = 2'b00;	 rom[3][21][1] = 2'b00;	 rom[3][22][1] = 2'b00;	 rom[3][23][1] = 2'b00;	 rom[3][24][1] = 2'b00;	 rom[3][25][1] = 2'b00;	 rom[3][26][1] = 2'b00;	 rom[3][27][1] = 2'b00;	 rom[3][28][1] = 2'b00;	 rom[3][29][1] = 2'b00;	 rom[3][30][1] = 2'b00;	 rom[3][31][1] = 2'b00;	 rom[3][32][1] = 2'b00;	 rom[3][33][1] = 2'b00;	 rom[3][34][1] = 2'b00;	 rom[3][35][1] = 2'b00;	 rom[3][36][1] = 2'b00;	 rom[3][37][1] = 2'b00;	 rom[3][38][1] = 2'b00;	 rom[3][39][1] = 2'b00;
 rom[3][0][2] = 2'b00;	 rom[3][1][2] = 2'b00;	 rom[3][2][2] = 2'b00;	 rom[3][3][2] = 2'b00;	 rom[3][4][2] = 2'b00;	 rom[3][5][2] = 2'b00;	 rom[3][6][2] = 2'b00;	 rom[3][7][2] = 2'b00;	 rom[3][8][2] = 2'b00;	 rom[3][9][2] = 2'b00;	 rom[3][10][2] = 2'b00;	 rom[3][11][2] = 2'b10;	 rom[3][12][2] = 2'b10;	 rom[3][13][2] = 2'b10;	 rom[3][14][2] = 2'b10;	 rom[3][15][2] = 2'b10;	 rom[3][16][2] = 2'b10;	 rom[3][17][2] = 2'b10;	 rom[3][18][2] = 2'b10;	 rom[3][19][2] = 2'b10;	 rom[3][20][2] = 2'b10;	 rom[3][21][2] = 2'b00;	 rom[3][22][2] = 2'b00;	 rom[3][23][2] = 2'b00;	 rom[3][24][2] = 2'b00;	 rom[3][25][2] = 2'b00;	 rom[3][26][2] = 2'b00;	 rom[3][27][2] = 2'b00;	 rom[3][28][2] = 2'b00;	 rom[3][29][2] = 2'b00;	 rom[3][30][2] = 2'b00;	 rom[3][31][2] = 2'b00;	 rom[3][32][2] = 2'b00;	 rom[3][33][2] = 2'b00;	 rom[3][34][2] = 2'b00;	 rom[3][35][2] = 2'b00;	 rom[3][36][2] = 2'b00;	 rom[3][37][2] = 2'b00;	 rom[3][38][2] = 2'b00;	 rom[3][39][2] = 2'b00;
 rom[3][0][3] = 2'b00;	 rom[3][1][3] = 2'b00;	 rom[3][2][3] = 2'b00;	 rom[3][3][3] = 2'b00;	 rom[3][4][3] = 2'b00;	 rom[3][5][3] = 2'b00;	 rom[3][6][3] = 2'b00;	 rom[3][7][3] = 2'b00;	 rom[3][8][3] = 2'b00;	 rom[3][9][3] = 2'b00;	 rom[3][10][3] = 2'b10;	 rom[3][11][3] = 2'b10;	 rom[3][12][3] = 2'b01;	 rom[3][13][3] = 2'b01;	 rom[3][14][3] = 2'b01;	 rom[3][15][3] = 2'b01;	 rom[3][16][3] = 2'b01;	 rom[3][17][3] = 2'b01;	 rom[3][18][3] = 2'b01;	 rom[3][19][3] = 2'b10;	 rom[3][20][3] = 2'b10;	 rom[3][21][3] = 2'b01;	 rom[3][22][3] = 2'b00;	 rom[3][23][3] = 2'b00;	 rom[3][24][3] = 2'b00;	 rom[3][25][3] = 2'b00;	 rom[3][26][3] = 2'b00;	 rom[3][27][3] = 2'b00;	 rom[3][28][3] = 2'b00;	 rom[3][29][3] = 2'b00;	 rom[3][30][3] = 2'b00;	 rom[3][31][3] = 2'b00;	 rom[3][32][3] = 2'b00;	 rom[3][33][3] = 2'b00;	 rom[3][34][3] = 2'b00;	 rom[3][35][3] = 2'b00;	 rom[3][36][3] = 2'b00;	 rom[3][37][3] = 2'b00;	 rom[3][38][3] = 2'b00;	 rom[3][39][3] = 2'b00;
 rom[3][0][4] = 2'b00;	 rom[3][1][4] = 2'b00;	 rom[3][2][4] = 2'b00;	 rom[3][3][4] = 2'b00;	 rom[3][4][4] = 2'b00;	 rom[3][5][4] = 2'b00;	 rom[3][6][4] = 2'b00;	 rom[3][7][4] = 2'b00;	 rom[3][8][4] = 2'b00;	 rom[3][9][4] = 2'b10;	 rom[3][10][4] = 2'b10;	 rom[3][11][4] = 2'b01;	 rom[3][12][4] = 2'b01;	 rom[3][13][4] = 2'b01;	 rom[3][14][4] = 2'b01;	 rom[3][15][4] = 2'b01;	 rom[3][16][4] = 2'b01;	 rom[3][17][4] = 2'b01;	 rom[3][18][4] = 2'b01;	 rom[3][19][4] = 2'b01;	 rom[3][20][4] = 2'b10;	 rom[3][21][4] = 2'b10;	 rom[3][22][4] = 2'b00;	 rom[3][23][4] = 2'b00;	 rom[3][24][4] = 2'b00;	 rom[3][25][4] = 2'b00;	 rom[3][26][4] = 2'b00;	 rom[3][27][4] = 2'b00;	 rom[3][28][4] = 2'b00;	 rom[3][29][4] = 2'b00;	 rom[3][30][4] = 2'b00;	 rom[3][31][4] = 2'b00;	 rom[3][32][4] = 2'b00;	 rom[3][33][4] = 2'b00;	 rom[3][34][4] = 2'b00;	 rom[3][35][4] = 2'b00;	 rom[3][36][4] = 2'b00;	 rom[3][37][4] = 2'b00;	 rom[3][38][4] = 2'b00;	 rom[3][39][4] = 2'b00;
 rom[3][0][5] = 2'b00;	 rom[3][1][5] = 2'b00;	 rom[3][2][5] = 2'b00;	 rom[3][3][5] = 2'b00;	 rom[3][4][5] = 2'b00;	 rom[3][5][5] = 2'b00;	 rom[3][6][5] = 2'b00;	 rom[3][7][5] = 2'b00;	 rom[3][8][5] = 2'b00;	 rom[3][9][5] = 2'b10;	 rom[3][10][5] = 2'b10;	 rom[3][11][5] = 2'b01;	 rom[3][12][5] = 2'b01;	 rom[3][13][5] = 2'b01;	 rom[3][14][5] = 2'b01;	 rom[3][15][5] = 2'b01;	 rom[3][16][5] = 2'b01;	 rom[3][17][5] = 2'b01;	 rom[3][18][5] = 2'b01;	 rom[3][19][5] = 2'b01;	 rom[3][20][5] = 2'b01;	 rom[3][21][5] = 2'b10;	 rom[3][22][5] = 2'b01;	 rom[3][23][5] = 2'b10;	 rom[3][24][5] = 2'b00;	 rom[3][25][5] = 2'b00;	 rom[3][26][5] = 2'b00;	 rom[3][27][5] = 2'b00;	 rom[3][28][5] = 2'b00;	 rom[3][29][5] = 2'b00;	 rom[3][30][5] = 2'b00;	 rom[3][31][5] = 2'b00;	 rom[3][32][5] = 2'b00;	 rom[3][33][5] = 2'b00;	 rom[3][34][5] = 2'b00;	 rom[3][35][5] = 2'b00;	 rom[3][36][5] = 2'b00;	 rom[3][37][5] = 2'b00;	 rom[3][38][5] = 2'b00;	 rom[3][39][5] = 2'b00;
 rom[3][0][6] = 2'b00;	 rom[3][1][6] = 2'b00;	 rom[3][2][6] = 2'b00;	 rom[3][3][6] = 2'b00;	 rom[3][4][6] = 2'b00;	 rom[3][5][6] = 2'b00;	 rom[3][6][6] = 2'b00;	 rom[3][7][6] = 2'b00;	 rom[3][8][6] = 2'b00;	 rom[3][9][6] = 2'b10;	 rom[3][10][6] = 2'b10;	 rom[3][11][6] = 2'b01;	 rom[3][12][6] = 2'b01;	 rom[3][13][6] = 2'b10;	 rom[3][14][6] = 2'b10;	 rom[3][15][6] = 2'b10;	 rom[3][16][6] = 2'b10;	 rom[3][17][6] = 2'b10;	 rom[3][18][6] = 2'b10;	 rom[3][19][6] = 2'b10;	 rom[3][20][6] = 2'b10;	 rom[3][21][6] = 2'b10;	 rom[3][22][6] = 2'b10;	 rom[3][23][6] = 2'b00;	 rom[3][24][6] = 2'b00;	 rom[3][25][6] = 2'b00;	 rom[3][26][6] = 2'b00;	 rom[3][27][6] = 2'b00;	 rom[3][28][6] = 2'b00;	 rom[3][29][6] = 2'b00;	 rom[3][30][6] = 2'b00;	 rom[3][31][6] = 2'b00;	 rom[3][32][6] = 2'b00;	 rom[3][33][6] = 2'b00;	 rom[3][34][6] = 2'b00;	 rom[3][35][6] = 2'b00;	 rom[3][36][6] = 2'b00;	 rom[3][37][6] = 2'b00;	 rom[3][38][6] = 2'b00;	 rom[3][39][6] = 2'b00;
 rom[3][0][7] = 2'b00;	 rom[3][1][7] = 2'b00;	 rom[3][2][7] = 2'b00;	 rom[3][3][7] = 2'b00;	 rom[3][4][7] = 2'b00;	 rom[3][5][7] = 2'b00;	 rom[3][6][7] = 2'b00;	 rom[3][7][7] = 2'b00;	 rom[3][8][7] = 2'b00;	 rom[3][9][7] = 2'b10;	 rom[3][10][7] = 2'b10;	 rom[3][11][7] = 2'b01;	 rom[3][12][7] = 2'b10;	 rom[3][13][7] = 2'b10;	 rom[3][14][7] = 2'b10;	 rom[3][15][7] = 2'b10;	 rom[3][16][7] = 2'b10;	 rom[3][17][7] = 2'b10;	 rom[3][18][7] = 2'b10;	 rom[3][19][7] = 2'b10;	 rom[3][20][7] = 2'b10;	 rom[3][21][7] = 2'b10;	 rom[3][22][7] = 2'b10;	 rom[3][23][7] = 2'b00;	 rom[3][24][7] = 2'b10;	 rom[3][25][7] = 2'b10;	 rom[3][26][7] = 2'b10;	 rom[3][27][7] = 2'b10;	 rom[3][28][7] = 2'b10;	 rom[3][29][7] = 2'b10;	 rom[3][30][7] = 2'b10;	 rom[3][31][7] = 2'b00;	 rom[3][32][7] = 2'b00;	 rom[3][33][7] = 2'b00;	 rom[3][34][7] = 2'b00;	 rom[3][35][7] = 2'b00;	 rom[3][36][7] = 2'b00;	 rom[3][37][7] = 2'b00;	 rom[3][38][7] = 2'b00;	 rom[3][39][7] = 2'b00;
 rom[3][0][8] = 2'b00;	 rom[3][1][8] = 2'b00;	 rom[3][2][8] = 2'b00;	 rom[3][3][8] = 2'b00;	 rom[3][4][8] = 2'b00;	 rom[3][5][8] = 2'b00;	 rom[3][6][8] = 2'b10;	 rom[3][7][8] = 2'b10;	 rom[3][8][8] = 2'b10;	 rom[3][9][8] = 2'b10;	 rom[3][10][8] = 2'b10;	 rom[3][11][8] = 2'b10;	 rom[3][12][8] = 2'b10;	 rom[3][13][8] = 2'b10;	 rom[3][14][8] = 2'b01;	 rom[3][15][8] = 2'b01;	 rom[3][16][8] = 2'b01;	 rom[3][17][8] = 2'b01;	 rom[3][18][8] = 2'b01;	 rom[3][19][8] = 2'b01;	 rom[3][20][8] = 2'b10;	 rom[3][21][8] = 2'b10;	 rom[3][22][8] = 2'b10;	 rom[3][23][8] = 2'b10;	 rom[3][24][8] = 2'b10;	 rom[3][25][8] = 2'b11;	 rom[3][26][8] = 2'b11;	 rom[3][27][8] = 2'b11;	 rom[3][28][8] = 2'b11;	 rom[3][29][8] = 2'b11;	 rom[3][30][8] = 2'b10;	 rom[3][31][8] = 2'b10;	 rom[3][32][8] = 2'b00;	 rom[3][33][8] = 2'b00;	 rom[3][34][8] = 2'b00;	 rom[3][35][8] = 2'b00;	 rom[3][36][8] = 2'b00;	 rom[3][37][8] = 2'b00;	 rom[3][38][8] = 2'b00;	 rom[3][39][8] = 2'b00;
 rom[3][0][9] = 2'b00;	 rom[3][1][9] = 2'b00;	 rom[3][2][9] = 2'b00;	 rom[3][3][9] = 2'b00;	 rom[3][4][9] = 2'b10;	 rom[3][5][9] = 2'b10;	 rom[3][6][9] = 2'b10;	 rom[3][7][9] = 2'b10;	 rom[3][8][9] = 2'b10;	 rom[3][9][9] = 2'b10;	 rom[3][10][9] = 2'b10;	 rom[3][11][9] = 2'b10;	 rom[3][12][9] = 2'b10;	 rom[3][13][9] = 2'b01;	 rom[3][14][9] = 2'b01;	 rom[3][15][9] = 2'b01;	 rom[3][16][9] = 2'b01;	 rom[3][17][9] = 2'b01;	 rom[3][18][9] = 2'b01;	 rom[3][19][9] = 2'b01;	 rom[3][20][9] = 2'b01;	 rom[3][21][9] = 2'b01;	 rom[3][22][9] = 2'b01;	 rom[3][23][9] = 2'b10;	 rom[3][24][9] = 2'b10;	 rom[3][25][9] = 2'b10;	 rom[3][26][9] = 2'b11;	 rom[3][27][9] = 2'b11;	 rom[3][28][9] = 2'b11;	 rom[3][29][9] = 2'b11;	 rom[3][30][9] = 2'b11;	 rom[3][31][9] = 2'b10;	 rom[3][32][9] = 2'b10;	 rom[3][33][9] = 2'b00;	 rom[3][34][9] = 2'b00;	 rom[3][35][9] = 2'b00;	 rom[3][36][9] = 2'b00;	 rom[3][37][9] = 2'b00;	 rom[3][38][9] = 2'b00;	 rom[3][39][9] = 2'b00;
 rom[3][0][10] = 2'b00;	 rom[3][1][10] = 2'b00;	 rom[3][2][10] = 2'b10;	 rom[3][3][10] = 2'b10;	 rom[3][4][10] = 2'b10;	 rom[3][5][10] = 2'b10;	 rom[3][6][10] = 2'b10;	 rom[3][7][10] = 2'b10;	 rom[3][8][10] = 2'b10;	 rom[3][9][10] = 2'b10;	 rom[3][10][10] = 2'b10;	 rom[3][11][10] = 2'b10;	 rom[3][12][10] = 2'b01;	 rom[3][13][10] = 2'b01;	 rom[3][14][10] = 2'b01;	 rom[3][15][10] = 2'b01;	 rom[3][16][10] = 2'b01;	 rom[3][17][10] = 2'b01;	 rom[3][18][10] = 2'b01;	 rom[3][19][10] = 2'b01;	 rom[3][20][10] = 2'b01;	 rom[3][21][10] = 2'b01;	 rom[3][22][10] = 2'b01;	 rom[3][23][10] = 2'b01;	 rom[3][24][10] = 2'b10;	 rom[3][25][10] = 2'b10;	 rom[3][26][10] = 2'b10;	 rom[3][27][10] = 2'b11;	 rom[3][28][10] = 2'b11;	 rom[3][29][10] = 2'b11;	 rom[3][30][10] = 2'b11;	 rom[3][31][10] = 2'b11;	 rom[3][32][10] = 2'b10;	 rom[3][33][10] = 2'b00;	 rom[3][34][10] = 2'b00;	 rom[3][35][10] = 2'b00;	 rom[3][36][10] = 2'b00;	 rom[3][37][10] = 2'b00;	 rom[3][38][10] = 2'b00;	 rom[3][39][10] = 2'b00;
 rom[3][0][11] = 2'b00;	 rom[3][1][11] = 2'b00;	 rom[3][2][11] = 2'b10;	 rom[3][3][11] = 2'b11;	 rom[3][4][11] = 2'b11;	 rom[3][5][11] = 2'b11;	 rom[3][6][11] = 2'b10;	 rom[3][7][11] = 2'b10;	 rom[3][8][11] = 2'b10;	 rom[3][9][11] = 2'b10;	 rom[3][10][11] = 2'b10;	 rom[3][11][11] = 2'b01;	 rom[3][12][11] = 2'b01;	 rom[3][13][11] = 2'b01;	 rom[3][14][11] = 2'b01;	 rom[3][15][11] = 2'b01;	 rom[3][16][11] = 2'b01;	 rom[3][17][11] = 2'b01;	 rom[3][18][11] = 2'b01;	 rom[3][19][11] = 2'b01;	 rom[3][20][11] = 2'b01;	 rom[3][21][11] = 2'b01;	 rom[3][22][11] = 2'b01;	 rom[3][23][11] = 2'b01;	 rom[3][24][11] = 2'b01;	 rom[3][25][11] = 2'b10;	 rom[3][26][11] = 2'b10;	 rom[3][27][11] = 2'b11;	 rom[3][28][11] = 2'b11;	 rom[3][29][11] = 2'b11;	 rom[3][30][11] = 2'b11;	 rom[3][31][11] = 2'b11;	 rom[3][32][11] = 2'b10;	 rom[3][33][11] = 2'b00;	 rom[3][34][11] = 2'b00;	 rom[3][35][11] = 2'b00;	 rom[3][36][11] = 2'b00;	 rom[3][37][11] = 2'b00;	 rom[3][38][11] = 2'b00;	 rom[3][39][11] = 2'b00;
 rom[3][0][12] = 2'b00;	 rom[3][1][12] = 2'b00;	 rom[3][2][12] = 2'b10;	 rom[3][3][12] = 2'b11;	 rom[3][4][12] = 2'b11;	 rom[3][5][12] = 2'b11;	 rom[3][6][12] = 2'b11;	 rom[3][7][12] = 2'b10;	 rom[3][8][12] = 2'b10;	 rom[3][9][12] = 2'b10;	 rom[3][10][12] = 2'b01;	 rom[3][11][12] = 2'b01;	 rom[3][12][12] = 2'b01;	 rom[3][13][12] = 2'b01;	 rom[3][14][12] = 2'b01;	 rom[3][15][12] = 2'b01;	 rom[3][16][12] = 2'b01;	 rom[3][17][12] = 2'b01;	 rom[3][18][12] = 2'b01;	 rom[3][19][12] = 2'b01;	 rom[3][20][12] = 2'b01;	 rom[3][21][12] = 2'b01;	 rom[3][22][12] = 2'b01;	 rom[3][23][12] = 2'b01;	 rom[3][24][12] = 2'b01;	 rom[3][25][12] = 2'b01;	 rom[3][26][12] = 2'b10;	 rom[3][27][12] = 2'b10;	 rom[3][28][12] = 2'b10;	 rom[3][29][12] = 2'b11;	 rom[3][30][12] = 2'b11;	 rom[3][31][12] = 2'b11;	 rom[3][32][12] = 2'b10;	 rom[3][33][12] = 2'b00;	 rom[3][34][12] = 2'b00;	 rom[3][35][12] = 2'b00;	 rom[3][36][12] = 2'b00;	 rom[3][37][12] = 2'b00;	 rom[3][38][12] = 2'b00;	 rom[3][39][12] = 2'b00;
 rom[3][0][13] = 2'b00;	 rom[3][1][13] = 2'b00;	 rom[3][2][13] = 2'b10;	 rom[3][3][13] = 2'b11;	 rom[3][4][13] = 2'b11;	 rom[3][5][13] = 2'b11;	 rom[3][6][13] = 2'b11;	 rom[3][7][13] = 2'b11;	 rom[3][8][13] = 2'b11;	 rom[3][9][13] = 2'b10;	 rom[3][10][13] = 2'b01;	 rom[3][11][13] = 2'b01;	 rom[3][12][13] = 2'b01;	 rom[3][13][13] = 2'b01;	 rom[3][14][13] = 2'b01;	 rom[3][15][13] = 2'b01;	 rom[3][16][13] = 2'b01;	 rom[3][17][13] = 2'b01;	 rom[3][18][13] = 2'b01;	 rom[3][19][13] = 2'b01;	 rom[3][20][13] = 2'b01;	 rom[3][21][13] = 2'b01;	 rom[3][22][13] = 2'b01;	 rom[3][23][13] = 2'b01;	 rom[3][24][13] = 2'b01;	 rom[3][25][13] = 2'b01;	 rom[3][26][13] = 2'b01;	 rom[3][27][13] = 2'b10;	 rom[3][28][13] = 2'b10;	 rom[3][29][13] = 2'b11;	 rom[3][30][13] = 2'b11;	 rom[3][31][13] = 2'b11;	 rom[3][32][13] = 2'b10;	 rom[3][33][13] = 2'b00;	 rom[3][34][13] = 2'b00;	 rom[3][35][13] = 2'b00;	 rom[3][36][13] = 2'b00;	 rom[3][37][13] = 2'b00;	 rom[3][38][13] = 2'b00;	 rom[3][39][13] = 2'b00;
 rom[3][0][14] = 2'b00;	 rom[3][1][14] = 2'b00;	 rom[3][2][14] = 2'b10;	 rom[3][3][14] = 2'b11;	 rom[3][4][14] = 2'b11;	 rom[3][5][14] = 2'b11;	 rom[3][6][14] = 2'b11;	 rom[3][7][14] = 2'b11;	 rom[3][8][14] = 2'b11;	 rom[3][9][14] = 2'b10;	 rom[3][10][14] = 2'b01;	 rom[3][11][14] = 2'b01;	 rom[3][12][14] = 2'b01;	 rom[3][13][14] = 2'b01;	 rom[3][14][14] = 2'b01;	 rom[3][15][14] = 2'b01;	 rom[3][16][14] = 2'b01;	 rom[3][17][14] = 2'b01;	 rom[3][18][14] = 2'b01;	 rom[3][19][14] = 2'b01;	 rom[3][20][14] = 2'b01;	 rom[3][21][14] = 2'b01;	 rom[3][22][14] = 2'b01;	 rom[3][23][14] = 2'b01;	 rom[3][24][14] = 2'b01;	 rom[3][25][14] = 2'b01;	 rom[3][26][14] = 2'b01;	 rom[3][27][14] = 2'b01;	 rom[3][28][14] = 2'b10;	 rom[3][29][14] = 2'b10;	 rom[3][30][14] = 2'b11;	 rom[3][31][14] = 2'b10;	 rom[3][32][14] = 2'b10;	 rom[3][33][14] = 2'b00;	 rom[3][34][14] = 2'b00;	 rom[3][35][14] = 2'b00;	 rom[3][36][14] = 2'b00;	 rom[3][37][14] = 2'b00;	 rom[3][38][14] = 2'b00;	 rom[3][39][14] = 2'b00;
 rom[3][0][15] = 2'b00;	 rom[3][1][15] = 2'b00;	 rom[3][2][15] = 2'b10;	 rom[3][3][15] = 2'b11;	 rom[3][4][15] = 2'b11;	 rom[3][5][15] = 2'b11;	 rom[3][6][15] = 2'b10;	 rom[3][7][15] = 2'b10;	 rom[3][8][15] = 2'b10;	 rom[3][9][15] = 2'b10;	 rom[3][10][15] = 2'b01;	 rom[3][11][15] = 2'b01;	 rom[3][12][15] = 2'b01;	 rom[3][13][15] = 2'b01;	 rom[3][14][15] = 2'b01;	 rom[3][15][15] = 2'b01;	 rom[3][16][15] = 2'b01;	 rom[3][17][15] = 2'b01;	 rom[3][18][15] = 2'b01;	 rom[3][19][15] = 2'b01;	 rom[3][20][15] = 2'b01;	 rom[3][21][15] = 2'b01;	 rom[3][22][15] = 2'b01;	 rom[3][23][15] = 2'b01;	 rom[3][24][15] = 2'b01;	 rom[3][25][15] = 2'b01;	 rom[3][26][15] = 2'b01;	 rom[3][27][15] = 2'b01;	 rom[3][28][15] = 2'b10;	 rom[3][29][15] = 2'b10;	 rom[3][30][15] = 2'b10;	 rom[3][31][15] = 2'b10;	 rom[3][32][15] = 2'b00;	 rom[3][33][15] = 2'b00;	 rom[3][34][15] = 2'b00;	 rom[3][35][15] = 2'b00;	 rom[3][36][15] = 2'b00;	 rom[3][37][15] = 2'b00;	 rom[3][38][15] = 2'b00;	 rom[3][39][15] = 2'b00;
 rom[3][0][16] = 2'b00;	 rom[3][1][16] = 2'b00;	 rom[3][2][16] = 2'b10;	 rom[3][3][16] = 2'b11;	 rom[3][4][16] = 2'b11;	 rom[3][5][16] = 2'b11;	 rom[3][6][16] = 2'b10;	 rom[3][7][16] = 2'b10;	 rom[3][8][16] = 2'b10;	 rom[3][9][16] = 2'b01;	 rom[3][10][16] = 2'b01;	 rom[3][11][16] = 2'b01;	 rom[3][12][16] = 2'b01;	 rom[3][13][16] = 2'b01;	 rom[3][14][16] = 2'b01;	 rom[3][15][16] = 2'b01;	 rom[3][16][16] = 2'b01;	 rom[3][17][16] = 2'b01;	 rom[3][18][16] = 2'b01;	 rom[3][19][16] = 2'b01;	 rom[3][20][16] = 2'b01;	 rom[3][21][16] = 2'b01;	 rom[3][22][16] = 2'b01;	 rom[3][23][16] = 2'b01;	 rom[3][24][16] = 2'b01;	 rom[3][25][16] = 2'b01;	 rom[3][26][16] = 2'b01;	 rom[3][27][16] = 2'b01;	 rom[3][28][16] = 2'b10;	 rom[3][29][16] = 2'b10;	 rom[3][30][16] = 2'b10;	 rom[3][31][16] = 2'b00;	 rom[3][32][16] = 2'b00;	 rom[3][33][16] = 2'b00;	 rom[3][34][16] = 2'b00;	 rom[3][35][16] = 2'b00;	 rom[3][36][16] = 2'b00;	 rom[3][37][16] = 2'b00;	 rom[3][38][16] = 2'b00;	 rom[3][39][16] = 2'b00;
 rom[3][0][17] = 2'b00;	 rom[3][1][17] = 2'b00;	 rom[3][2][17] = 2'b10;	 rom[3][3][17] = 2'b11;	 rom[3][4][17] = 2'b10;	 rom[3][5][17] = 2'b11;	 rom[3][6][17] = 2'b10;	 rom[3][7][17] = 2'b10;	 rom[3][8][17] = 2'b10;	 rom[3][9][17] = 2'b01;	 rom[3][10][17] = 2'b01;	 rom[3][11][17] = 2'b01;	 rom[3][12][17] = 2'b01;	 rom[3][13][17] = 2'b01;	 rom[3][14][17] = 2'b01;	 rom[3][15][17] = 2'b01;	 rom[3][16][17] = 2'b01;	 rom[3][17][17] = 2'b01;	 rom[3][18][17] = 2'b01;	 rom[3][19][17] = 2'b01;	 rom[3][20][17] = 2'b01;	 rom[3][21][17] = 2'b01;	 rom[3][22][17] = 2'b01;	 rom[3][23][17] = 2'b01;	 rom[3][24][17] = 2'b01;	 rom[3][25][17] = 2'b01;	 rom[3][26][17] = 2'b01;	 rom[3][27][17] = 2'b01;	 rom[3][28][17] = 2'b10;	 rom[3][29][17] = 2'b10;	 rom[3][30][17] = 2'b00;	 rom[3][31][17] = 2'b00;	 rom[3][32][17] = 2'b00;	 rom[3][33][17] = 2'b00;	 rom[3][34][17] = 2'b00;	 rom[3][35][17] = 2'b00;	 rom[3][36][17] = 2'b00;	 rom[3][37][17] = 2'b00;	 rom[3][38][17] = 2'b00;	 rom[3][39][17] = 2'b00;
 rom[3][0][18] = 2'b00;	 rom[3][1][18] = 2'b00;	 rom[3][2][18] = 2'b10;	 rom[3][3][18] = 2'b11;	 rom[3][4][18] = 2'b10;	 rom[3][5][18] = 2'b11;	 rom[3][6][18] = 2'b10;	 rom[3][7][18] = 2'b10;	 rom[3][8][18] = 2'b10;	 rom[3][9][18] = 2'b01;	 rom[3][10][18] = 2'b01;	 rom[3][11][18] = 2'b01;	 rom[3][12][18] = 2'b01;	 rom[3][13][18] = 2'b01;	 rom[3][14][18] = 2'b01;	 rom[3][15][18] = 2'b01;	 rom[3][16][18] = 2'b01;	 rom[3][17][18] = 2'b01;	 rom[3][18][18] = 2'b01;	 rom[3][19][18] = 2'b01;	 rom[3][20][18] = 2'b01;	 rom[3][21][18] = 2'b01;	 rom[3][22][18] = 2'b01;	 rom[3][23][18] = 2'b01;	 rom[3][24][18] = 2'b01;	 rom[3][25][18] = 2'b01;	 rom[3][26][18] = 2'b01;	 rom[3][27][18] = 2'b01;	 rom[3][28][18] = 2'b10;	 rom[3][29][18] = 2'b10;	 rom[3][30][18] = 2'b10;	 rom[3][31][18] = 2'b10;	 rom[3][32][18] = 2'b10;	 rom[3][33][18] = 2'b00;	 rom[3][34][18] = 2'b00;	 rom[3][35][18] = 2'b00;	 rom[3][36][18] = 2'b00;	 rom[3][37][18] = 2'b00;	 rom[3][38][18] = 2'b00;	 rom[3][39][18] = 2'b00;
 rom[3][0][19] = 2'b00;	 rom[3][1][19] = 2'b00;	 rom[3][2][19] = 2'b10;	 rom[3][3][19] = 2'b11;	 rom[3][4][19] = 2'b10;	 rom[3][5][19] = 2'b11;	 rom[3][6][19] = 2'b10;	 rom[3][7][19] = 2'b10;	 rom[3][8][19] = 2'b10;	 rom[3][9][19] = 2'b01;	 rom[3][10][19] = 2'b01;	 rom[3][11][19] = 2'b01;	 rom[3][12][19] = 2'b01;	 rom[3][13][19] = 2'b01;	 rom[3][14][19] = 2'b01;	 rom[3][15][19] = 2'b01;	 rom[3][16][19] = 2'b01;	 rom[3][17][19] = 2'b01;	 rom[3][18][19] = 2'b01;	 rom[3][19][19] = 2'b01;	 rom[3][20][19] = 2'b01;	 rom[3][21][19] = 2'b01;	 rom[3][22][19] = 2'b01;	 rom[3][23][19] = 2'b01;	 rom[3][24][19] = 2'b01;	 rom[3][25][19] = 2'b01;	 rom[3][26][19] = 2'b01;	 rom[3][27][19] = 2'b01;	 rom[3][28][19] = 2'b10;	 rom[3][29][19] = 2'b10;	 rom[3][30][19] = 2'b11;	 rom[3][31][19] = 2'b11;	 rom[3][32][19] = 2'b10;	 rom[3][33][19] = 2'b10;	 rom[3][34][19] = 2'b00;	 rom[3][35][19] = 2'b00;	 rom[3][36][19] = 2'b00;	 rom[3][37][19] = 2'b00;	 rom[3][38][19] = 2'b00;	 rom[3][39][19] = 2'b00;
 rom[3][0][20] = 2'b00;	 rom[3][1][20] = 2'b00;	 rom[3][2][20] = 2'b10;	 rom[3][3][20] = 2'b11;	 rom[3][4][20] = 2'b10;	 rom[3][5][20] = 2'b11;	 rom[3][6][20] = 2'b10;	 rom[3][7][20] = 2'b10;	 rom[3][8][20] = 2'b10;	 rom[3][9][20] = 2'b01;	 rom[3][10][20] = 2'b01;	 rom[3][11][20] = 2'b01;	 rom[3][12][20] = 2'b01;	 rom[3][13][20] = 2'b01;	 rom[3][14][20] = 2'b01;	 rom[3][15][20] = 2'b01;	 rom[3][16][20] = 2'b01;	 rom[3][17][20] = 2'b01;	 rom[3][18][20] = 2'b01;	 rom[3][19][20] = 2'b01;	 rom[3][20][20] = 2'b01;	 rom[3][21][20] = 2'b01;	 rom[3][22][20] = 2'b01;	 rom[3][23][20] = 2'b01;	 rom[3][24][20] = 2'b01;	 rom[3][25][20] = 2'b01;	 rom[3][26][20] = 2'b01;	 rom[3][27][20] = 2'b01;	 rom[3][28][20] = 2'b10;	 rom[3][29][20] = 2'b10;	 rom[3][30][20] = 2'b11;	 rom[3][31][20] = 2'b11;	 rom[3][32][20] = 2'b11;	 rom[3][33][20] = 2'b10;	 rom[3][34][20] = 2'b00;	 rom[3][35][20] = 2'b00;	 rom[3][36][20] = 2'b00;	 rom[3][37][20] = 2'b00;	 rom[3][38][20] = 2'b00;	 rom[3][39][20] = 2'b00;
 rom[3][0][21] = 2'b00;	 rom[3][1][21] = 2'b00;	 rom[3][2][21] = 2'b10;	 rom[3][3][21] = 2'b11;	 rom[3][4][21] = 2'b10;	 rom[3][5][21] = 2'b11;	 rom[3][6][21] = 2'b10;	 rom[3][7][21] = 2'b10;	 rom[3][8][21] = 2'b10;	 rom[3][9][21] = 2'b01;	 rom[3][10][21] = 2'b01;	 rom[3][11][21] = 2'b01;	 rom[3][12][21] = 2'b01;	 rom[3][13][21] = 2'b01;	 rom[3][14][21] = 2'b01;	 rom[3][15][21] = 2'b01;	 rom[3][16][21] = 2'b01;	 rom[3][17][21] = 2'b01;	 rom[3][18][21] = 2'b01;	 rom[3][19][21] = 2'b01;	 rom[3][20][21] = 2'b01;	 rom[3][21][21] = 2'b01;	 rom[3][22][21] = 2'b01;	 rom[3][23][21] = 2'b01;	 rom[3][24][21] = 2'b01;	 rom[3][25][21] = 2'b01;	 rom[3][26][21] = 2'b01;	 rom[3][27][21] = 2'b01;	 rom[3][28][21] = 2'b10;	 rom[3][29][21] = 2'b10;	 rom[3][30][21] = 2'b11;	 rom[3][31][21] = 2'b11;	 rom[3][32][21] = 2'b11;	 rom[3][33][21] = 2'b10;	 rom[3][34][21] = 2'b00;	 rom[3][35][21] = 2'b00;	 rom[3][36][21] = 2'b00;	 rom[3][37][21] = 2'b00;	 rom[3][38][21] = 2'b00;	 rom[3][39][21] = 2'b00;
 rom[3][0][22] = 2'b00;	 rom[3][1][22] = 2'b00;	 rom[3][2][22] = 2'b10;	 rom[3][3][22] = 2'b11;	 rom[3][4][22] = 2'b10;	 rom[3][5][22] = 2'b11;	 rom[3][6][22] = 2'b10;	 rom[3][7][22] = 2'b10;	 rom[3][8][22] = 2'b10;	 rom[3][9][22] = 2'b01;	 rom[3][10][22] = 2'b01;	 rom[3][11][22] = 2'b01;	 rom[3][12][22] = 2'b01;	 rom[3][13][22] = 2'b01;	 rom[3][14][22] = 2'b01;	 rom[3][15][22] = 2'b01;	 rom[3][16][22] = 2'b01;	 rom[3][17][22] = 2'b01;	 rom[3][18][22] = 2'b01;	 rom[3][19][22] = 2'b01;	 rom[3][20][22] = 2'b01;	 rom[3][21][22] = 2'b01;	 rom[3][22][22] = 2'b01;	 rom[3][23][22] = 2'b01;	 rom[3][24][22] = 2'b01;	 rom[3][25][22] = 2'b01;	 rom[3][26][22] = 2'b01;	 rom[3][27][22] = 2'b01;	 rom[3][28][22] = 2'b10;	 rom[3][29][22] = 2'b10;	 rom[3][30][22] = 2'b11;	 rom[3][31][22] = 2'b11;	 rom[3][32][22] = 2'b11;	 rom[3][33][22] = 2'b10;	 rom[3][34][22] = 2'b00;	 rom[3][35][22] = 2'b00;	 rom[3][36][22] = 2'b00;	 rom[3][37][22] = 2'b00;	 rom[3][38][22] = 2'b00;	 rom[3][39][22] = 2'b00;
 rom[3][0][23] = 2'b00;	 rom[3][1][23] = 2'b00;	 rom[3][2][23] = 2'b10;	 rom[3][3][23] = 2'b11;	 rom[3][4][23] = 2'b11;	 rom[3][5][23] = 2'b11;	 rom[3][6][23] = 2'b10;	 rom[3][7][23] = 2'b10;	 rom[3][8][23] = 2'b10;	 rom[3][9][23] = 2'b01;	 rom[3][10][23] = 2'b01;	 rom[3][11][23] = 2'b01;	 rom[3][12][23] = 2'b01;	 rom[3][13][23] = 2'b01;	 rom[3][14][23] = 2'b01;	 rom[3][15][23] = 2'b01;	 rom[3][16][23] = 2'b01;	 rom[3][17][23] = 2'b01;	 rom[3][18][23] = 2'b01;	 rom[3][19][23] = 2'b01;	 rom[3][20][23] = 2'b01;	 rom[3][21][23] = 2'b01;	 rom[3][22][23] = 2'b01;	 rom[3][23][23] = 2'b01;	 rom[3][24][23] = 2'b01;	 rom[3][25][23] = 2'b01;	 rom[3][26][23] = 2'b01;	 rom[3][27][23] = 2'b01;	 rom[3][28][23] = 2'b10;	 rom[3][29][23] = 2'b10;	 rom[3][30][23] = 2'b11;	 rom[3][31][23] = 2'b11;	 rom[3][32][23] = 2'b11;	 rom[3][33][23] = 2'b10;	 rom[3][34][23] = 2'b00;	 rom[3][35][23] = 2'b00;	 rom[3][36][23] = 2'b00;	 rom[3][37][23] = 2'b00;	 rom[3][38][23] = 2'b00;	 rom[3][39][23] = 2'b00;
 rom[3][0][24] = 2'b00;	 rom[3][1][24] = 2'b00;	 rom[3][2][24] = 2'b10;	 rom[3][3][24] = 2'b11;	 rom[3][4][24] = 2'b11;	 rom[3][5][24] = 2'b11;	 rom[3][6][24] = 2'b10;	 rom[3][7][24] = 2'b10;	 rom[3][8][24] = 2'b10;	 rom[3][9][24] = 2'b10;	 rom[3][10][24] = 2'b01;	 rom[3][11][24] = 2'b01;	 rom[3][12][24] = 2'b01;	 rom[3][13][24] = 2'b01;	 rom[3][14][24] = 2'b01;	 rom[3][15][24] = 2'b01;	 rom[3][16][24] = 2'b01;	 rom[3][17][24] = 2'b01;	 rom[3][18][24] = 2'b01;	 rom[3][19][24] = 2'b01;	 rom[3][20][24] = 2'b01;	 rom[3][21][24] = 2'b01;	 rom[3][22][24] = 2'b01;	 rom[3][23][24] = 2'b01;	 rom[3][24][24] = 2'b01;	 rom[3][25][24] = 2'b01;	 rom[3][26][24] = 2'b01;	 rom[3][27][24] = 2'b01;	 rom[3][28][24] = 2'b10;	 rom[3][29][24] = 2'b10;	 rom[3][30][24] = 2'b11;	 rom[3][31][24] = 2'b11;	 rom[3][32][24] = 2'b10;	 rom[3][33][24] = 2'b10;	 rom[3][34][24] = 2'b00;	 rom[3][35][24] = 2'b00;	 rom[3][36][24] = 2'b00;	 rom[3][37][24] = 2'b00;	 rom[3][38][24] = 2'b00;	 rom[3][39][24] = 2'b00;
 rom[3][0][25] = 2'b00;	 rom[3][1][25] = 2'b00;	 rom[3][2][25] = 2'b10;	 rom[3][3][25] = 2'b11;	 rom[3][4][25] = 2'b11;	 rom[3][5][25] = 2'b11;	 rom[3][6][25] = 2'b11;	 rom[3][7][25] = 2'b11;	 rom[3][8][25] = 2'b11;	 rom[3][9][25] = 2'b10;	 rom[3][10][25] = 2'b01;	 rom[3][11][25] = 2'b01;	 rom[3][12][25] = 2'b01;	 rom[3][13][25] = 2'b01;	 rom[3][14][25] = 2'b01;	 rom[3][15][25] = 2'b01;	 rom[3][16][25] = 2'b01;	 rom[3][17][25] = 2'b01;	 rom[3][18][25] = 2'b01;	 rom[3][19][25] = 2'b01;	 rom[3][20][25] = 2'b01;	 rom[3][21][25] = 2'b01;	 rom[3][22][25] = 2'b01;	 rom[3][23][25] = 2'b01;	 rom[3][24][25] = 2'b01;	 rom[3][25][25] = 2'b01;	 rom[3][26][25] = 2'b01;	 rom[3][27][25] = 2'b01;	 rom[3][28][25] = 2'b10;	 rom[3][29][25] = 2'b10;	 rom[3][30][25] = 2'b11;	 rom[3][31][25] = 2'b10;	 rom[3][32][25] = 2'b10;	 rom[3][33][25] = 2'b00;	 rom[3][34][25] = 2'b00;	 rom[3][35][25] = 2'b00;	 rom[3][36][25] = 2'b00;	 rom[3][37][25] = 2'b00;	 rom[3][38][25] = 2'b00;	 rom[3][39][25] = 2'b00;
 rom[3][0][26] = 2'b00;	 rom[3][1][26] = 2'b00;	 rom[3][2][26] = 2'b10;	 rom[3][3][26] = 2'b11;	 rom[3][4][26] = 2'b11;	 rom[3][5][26] = 2'b11;	 rom[3][6][26] = 2'b11;	 rom[3][7][26] = 2'b11;	 rom[3][8][26] = 2'b11;	 rom[3][9][26] = 2'b10;	 rom[3][10][26] = 2'b01;	 rom[3][11][26] = 2'b01;	 rom[3][12][26] = 2'b01;	 rom[3][13][26] = 2'b01;	 rom[3][14][26] = 2'b01;	 rom[3][15][26] = 2'b01;	 rom[3][16][26] = 2'b01;	 rom[3][17][26] = 2'b01;	 rom[3][18][26] = 2'b01;	 rom[3][19][26] = 2'b01;	 rom[3][20][26] = 2'b01;	 rom[3][21][26] = 2'b01;	 rom[3][22][26] = 2'b01;	 rom[3][23][26] = 2'b01;	 rom[3][24][26] = 2'b01;	 rom[3][25][26] = 2'b01;	 rom[3][26][26] = 2'b01;	 rom[3][27][26] = 2'b10;	 rom[3][28][26] = 2'b10;	 rom[3][29][26] = 2'b10;	 rom[3][30][26] = 2'b10;	 rom[3][31][26] = 2'b10;	 rom[3][32][26] = 2'b00;	 rom[3][33][26] = 2'b00;	 rom[3][34][26] = 2'b00;	 rom[3][35][26] = 2'b00;	 rom[3][36][26] = 2'b00;	 rom[3][37][26] = 2'b00;	 rom[3][38][26] = 2'b00;	 rom[3][39][26] = 2'b00;
 rom[3][0][27] = 2'b00;	 rom[3][1][27] = 2'b00;	 rom[3][2][27] = 2'b10;	 rom[3][3][27] = 2'b11;	 rom[3][4][27] = 2'b11;	 rom[3][5][27] = 2'b11;	 rom[3][6][27] = 2'b11;	 rom[3][7][27] = 2'b10;	 rom[3][8][27] = 2'b10;	 rom[3][9][27] = 2'b10;	 rom[3][10][27] = 2'b01;	 rom[3][11][27] = 2'b01;	 rom[3][12][27] = 2'b01;	 rom[3][13][27] = 2'b01;	 rom[3][14][27] = 2'b01;	 rom[3][15][27] = 2'b01;	 rom[3][16][27] = 2'b01;	 rom[3][17][27] = 2'b01;	 rom[3][18][27] = 2'b01;	 rom[3][19][27] = 2'b01;	 rom[3][20][27] = 2'b01;	 rom[3][21][27] = 2'b01;	 rom[3][22][27] = 2'b01;	 rom[3][23][27] = 2'b01;	 rom[3][24][27] = 2'b01;	 rom[3][25][27] = 2'b01;	 rom[3][26][27] = 2'b10;	 rom[3][27][27] = 2'b10;	 rom[3][28][27] = 2'b10;	 rom[3][29][27] = 2'b00;	 rom[3][30][27] = 2'b00;	 rom[3][31][27] = 2'b00;	 rom[3][32][27] = 2'b00;	 rom[3][33][27] = 2'b00;	 rom[3][34][27] = 2'b00;	 rom[3][35][27] = 2'b00;	 rom[3][36][27] = 2'b00;	 rom[3][37][27] = 2'b00;	 rom[3][38][27] = 2'b00;	 rom[3][39][27] = 2'b00;
 rom[3][0][28] = 2'b00;	 rom[3][1][28] = 2'b00;	 rom[3][2][28] = 2'b10;	 rom[3][3][28] = 2'b11;	 rom[3][4][28] = 2'b11;	 rom[3][5][28] = 2'b11;	 rom[3][6][28] = 2'b10;	 rom[3][7][28] = 2'b10;	 rom[3][8][28] = 2'b10;	 rom[3][9][28] = 2'b10;	 rom[3][10][28] = 2'b10;	 rom[3][11][28] = 2'b01;	 rom[3][12][28] = 2'b01;	 rom[3][13][28] = 2'b01;	 rom[3][14][28] = 2'b01;	 rom[3][15][28] = 2'b01;	 rom[3][16][28] = 2'b01;	 rom[3][17][28] = 2'b01;	 rom[3][18][28] = 2'b01;	 rom[3][19][28] = 2'b01;	 rom[3][20][28] = 2'b01;	 rom[3][21][28] = 2'b01;	 rom[3][22][28] = 2'b01;	 rom[3][23][28] = 2'b01;	 rom[3][24][28] = 2'b01;	 rom[3][25][28] = 2'b10;	 rom[3][26][28] = 2'b10;	 rom[3][27][28] = 2'b00;	 rom[3][28][28] = 2'b00;	 rom[3][29][28] = 2'b00;	 rom[3][30][28] = 2'b00;	 rom[3][31][28] = 2'b00;	 rom[3][32][28] = 2'b00;	 rom[3][33][28] = 2'b00;	 rom[3][34][28] = 2'b00;	 rom[3][35][28] = 2'b00;	 rom[3][36][28] = 2'b00;	 rom[3][37][28] = 2'b00;	 rom[3][38][28] = 2'b10;	 rom[3][39][28] = 2'b10;
 rom[3][0][29] = 2'b00;	 rom[3][1][29] = 2'b00;	 rom[3][2][29] = 2'b10;	 rom[3][3][29] = 2'b10;	 rom[3][4][29] = 2'b10;	 rom[3][5][29] = 2'b10;	 rom[3][6][29] = 2'b10;	 rom[3][7][29] = 2'b10;	 rom[3][8][29] = 2'b10;	 rom[3][9][29] = 2'b10;	 rom[3][10][29] = 2'b10;	 rom[3][11][29] = 2'b10;	 rom[3][12][29] = 2'b01;	 rom[3][13][29] = 2'b01;	 rom[3][14][29] = 2'b01;	 rom[3][15][29] = 2'b01;	 rom[3][16][29] = 2'b01;	 rom[3][17][29] = 2'b01;	 rom[3][18][29] = 2'b01;	 rom[3][19][29] = 2'b01;	 rom[3][20][29] = 2'b01;	 rom[3][21][29] = 2'b01;	 rom[3][22][29] = 2'b01;	 rom[3][23][29] = 2'b01;	 rom[3][24][29] = 2'b10;	 rom[3][25][29] = 2'b10;	 rom[3][26][29] = 2'b10;	 rom[3][27][29] = 2'b10;	 rom[3][28][29] = 2'b10;	 rom[3][29][29] = 2'b10;	 rom[3][30][29] = 2'b10;	 rom[3][31][29] = 2'b10;	 rom[3][32][29] = 2'b10;	 rom[3][33][29] = 2'b10;	 rom[3][34][29] = 2'b10;	 rom[3][35][29] = 2'b10;	 rom[3][36][29] = 2'b10;	 rom[3][37][29] = 2'b10;	 rom[3][38][29] = 2'b10;	 rom[3][39][29] = 2'b10;
 rom[3][0][30] = 2'b00;	 rom[3][1][30] = 2'b00;	 rom[3][2][30] = 2'b00;	 rom[3][3][30] = 2'b00;	 rom[3][4][30] = 2'b10;	 rom[3][5][30] = 2'b10;	 rom[3][6][30] = 2'b10;	 rom[3][7][30] = 2'b10;	 rom[3][8][30] = 2'b10;	 rom[3][9][30] = 2'b10;	 rom[3][10][30] = 2'b10;	 rom[3][11][30] = 2'b10;	 rom[3][12][30] = 2'b10;	 rom[3][13][30] = 2'b01;	 rom[3][14][30] = 2'b01;	 rom[3][15][30] = 2'b01;	 rom[3][16][30] = 2'b01;	 rom[3][17][30] = 2'b01;	 rom[3][18][30] = 2'b01;	 rom[3][19][30] = 2'b01;	 rom[3][20][30] = 2'b01;	 rom[3][21][30] = 2'b01;	 rom[3][22][30] = 2'b01;	 rom[3][23][30] = 2'b10;	 rom[3][24][30] = 2'b10;	 rom[3][25][30] = 2'b11;	 rom[3][26][30] = 2'b11;	 rom[3][27][30] = 2'b11;	 rom[3][28][30] = 2'b11;	 rom[3][29][30] = 2'b11;	 rom[3][30][30] = 2'b11;	 rom[3][31][30] = 2'b11;	 rom[3][32][30] = 2'b11;	 rom[3][33][30] = 2'b11;	 rom[3][34][30] = 2'b11;	 rom[3][35][30] = 2'b11;	 rom[3][36][30] = 2'b11;	 rom[3][37][30] = 2'b11;	 rom[3][38][30] = 2'b11;	 rom[3][39][30] = 2'b10;
 rom[3][0][31] = 2'b00;	 rom[3][1][31] = 2'b00;	 rom[3][2][31] = 2'b00;	 rom[3][3][31] = 2'b00;	 rom[3][4][31] = 2'b00;	 rom[3][5][31] = 2'b00;	 rom[3][6][31] = 2'b10;	 rom[3][7][31] = 2'b10;	 rom[3][8][31] = 2'b10;	 rom[3][9][31] = 2'b10;	 rom[3][10][31] = 2'b10;	 rom[3][11][31] = 2'b10;	 rom[3][12][31] = 2'b10;	 rom[3][13][31] = 2'b10;	 rom[3][14][31] = 2'b10;	 rom[3][15][31] = 2'b01;	 rom[3][16][31] = 2'b01;	 rom[3][17][31] = 2'b10;	 rom[3][18][31] = 2'b01;	 rom[3][19][31] = 2'b01;	 rom[3][20][31] = 2'b10;	 rom[3][21][31] = 2'b10;	 rom[3][22][31] = 2'b10;	 rom[3][23][31] = 2'b10;	 rom[3][24][31] = 2'b11;	 rom[3][25][31] = 2'b11;	 rom[3][26][31] = 2'b11;	 rom[3][27][31] = 2'b11;	 rom[3][28][31] = 2'b11;	 rom[3][29][31] = 2'b11;	 rom[3][30][31] = 2'b11;	 rom[3][31][31] = 2'b11;	 rom[3][32][31] = 2'b11;	 rom[3][33][31] = 2'b11;	 rom[3][34][31] = 2'b11;	 rom[3][35][31] = 2'b11;	 rom[3][36][31] = 2'b11;	 rom[3][37][31] = 2'b11;	 rom[3][38][31] = 2'b11;	 rom[3][39][31] = 2'b10;
 rom[3][0][32] = 2'b00;	 rom[3][1][32] = 2'b00;	 rom[3][2][32] = 2'b00;	 rom[3][3][32] = 2'b00;	 rom[3][4][32] = 2'b00;	 rom[3][5][32] = 2'b00;	 rom[3][6][32] = 2'b00;	 rom[3][7][32] = 2'b00;	 rom[3][8][32] = 2'b00;	 rom[3][9][32] = 2'b10;	 rom[3][10][32] = 2'b10;	 rom[3][11][32] = 2'b01;	 rom[3][12][32] = 2'b10;	 rom[3][13][32] = 2'b10;	 rom[3][14][32] = 2'b10;	 rom[3][15][32] = 2'b10;	 rom[3][16][32] = 2'b10;	 rom[3][17][32] = 2'b10;	 rom[3][18][32] = 2'b10;	 rom[3][19][32] = 2'b10;	 rom[3][20][32] = 2'b10;	 rom[3][21][32] = 2'b10;	 rom[3][22][32] = 2'b10;	 rom[3][23][32] = 2'b10;	 rom[3][24][32] = 2'b10;	 rom[3][25][32] = 2'b10;	 rom[3][26][32] = 2'b10;	 rom[3][27][32] = 2'b10;	 rom[3][28][32] = 2'b10;	 rom[3][29][32] = 2'b10;	 rom[3][30][32] = 2'b10;	 rom[3][31][32] = 2'b10;	 rom[3][32][32] = 2'b10;	 rom[3][33][32] = 2'b10;	 rom[3][34][32] = 2'b10;	 rom[3][35][32] = 2'b10;	 rom[3][36][32] = 2'b10;	 rom[3][37][32] = 2'b10;	 rom[3][38][32] = 2'b10;	 rom[3][39][32] = 2'b10;
 rom[3][0][33] = 2'b00;	 rom[3][1][33] = 2'b00;	 rom[3][2][33] = 2'b00;	 rom[3][3][33] = 2'b00;	 rom[3][4][33] = 2'b00;	 rom[3][5][33] = 2'b00;	 rom[3][6][33] = 2'b00;	 rom[3][7][33] = 2'b00;	 rom[3][8][33] = 2'b00;	 rom[3][9][33] = 2'b10;	 rom[3][10][33] = 2'b10;	 rom[3][11][33] = 2'b01;	 rom[3][12][33] = 2'b01;	 rom[3][13][33] = 2'b10;	 rom[3][14][33] = 2'b10;	 rom[3][15][33] = 2'b10;	 rom[3][16][33] = 2'b10;	 rom[3][17][33] = 2'b10;	 rom[3][18][33] = 2'b10;	 rom[3][19][33] = 2'b10;	 rom[3][20][33] = 2'b10;	 rom[3][21][33] = 2'b10;	 rom[3][22][33] = 2'b10;	 rom[3][23][33] = 2'b10;	 rom[3][24][33] = 2'b10;	 rom[3][25][33] = 2'b10;	 rom[3][26][33] = 2'b01;	 rom[3][27][33] = 2'b01;	 rom[3][28][33] = 2'b01;	 rom[3][29][33] = 2'b01;	 rom[3][30][33] = 2'b10;	 rom[3][31][33] = 2'b10;	 rom[3][32][33] = 2'b00;	 rom[3][33][33] = 2'b00;	 rom[3][34][33] = 2'b00;	 rom[3][35][33] = 2'b00;	 rom[3][36][33] = 2'b00;	 rom[3][37][33] = 2'b00;	 rom[3][38][33] = 2'b00;	 rom[3][39][33] = 2'b00;
 rom[3][0][34] = 2'b00;	 rom[3][1][34] = 2'b00;	 rom[3][2][34] = 2'b00;	 rom[3][3][34] = 2'b00;	 rom[3][4][34] = 2'b00;	 rom[3][5][34] = 2'b00;	 rom[3][6][34] = 2'b00;	 rom[3][7][34] = 2'b00;	 rom[3][8][34] = 2'b00;	 rom[3][9][34] = 2'b10;	 rom[3][10][34] = 2'b10;	 rom[3][11][34] = 2'b01;	 rom[3][12][34] = 2'b01;	 rom[3][13][34] = 2'b01;	 rom[3][14][34] = 2'b01;	 rom[3][15][34] = 2'b01;	 rom[3][16][34] = 2'b01;	 rom[3][17][34] = 2'b01;	 rom[3][18][34] = 2'b01;	 rom[3][19][34] = 2'b01;	 rom[3][20][34] = 2'b01;	 rom[3][21][34] = 2'b01;	 rom[3][22][34] = 2'b01;	 rom[3][23][34] = 2'b01;	 rom[3][24][34] = 2'b01;	 rom[3][25][34] = 2'b01;	 rom[3][26][34] = 2'b01;	 rom[3][27][34] = 2'b01;	 rom[3][28][34] = 2'b10;	 rom[3][29][34] = 2'b10;	 rom[3][30][34] = 2'b10;	 rom[3][31][34] = 2'b00;	 rom[3][32][34] = 2'b00;	 rom[3][33][34] = 2'b00;	 rom[3][34][34] = 2'b00;	 rom[3][35][34] = 2'b00;	 rom[3][36][34] = 2'b00;	 rom[3][37][34] = 2'b00;	 rom[3][38][34] = 2'b00;	 rom[3][39][34] = 2'b00;
 rom[3][0][35] = 2'b00;	 rom[3][1][35] = 2'b00;	 rom[3][2][35] = 2'b00;	 rom[3][3][35] = 2'b00;	 rom[3][4][35] = 2'b00;	 rom[3][5][35] = 2'b00;	 rom[3][6][35] = 2'b00;	 rom[3][7][35] = 2'b01;	 rom[3][8][35] = 2'b01;	 rom[3][9][35] = 2'b10;	 rom[3][10][35] = 2'b10;	 rom[3][11][35] = 2'b01;	 rom[3][12][35] = 2'b01;	 rom[3][13][35] = 2'b01;	 rom[3][14][35] = 2'b01;	 rom[3][15][35] = 2'b01;	 rom[3][16][35] = 2'b01;	 rom[3][17][35] = 2'b01;	 rom[3][18][35] = 2'b01;	 rom[3][19][35] = 2'b01;	 rom[3][20][35] = 2'b01;	 rom[3][21][35] = 2'b01;	 rom[3][22][35] = 2'b01;	 rom[3][23][35] = 2'b01;	 rom[3][24][35] = 2'b01;	 rom[3][25][35] = 2'b01;	 rom[3][26][35] = 2'b01;	 rom[3][27][35] = 2'b10;	 rom[3][28][35] = 2'b10;	 rom[3][29][35] = 2'b00;	 rom[3][30][35] = 2'b00;	 rom[3][31][35] = 2'b00;	 rom[3][32][35] = 2'b00;	 rom[3][33][35] = 2'b00;	 rom[3][34][35] = 2'b00;	 rom[3][35][35] = 2'b00;	 rom[3][36][35] = 2'b00;	 rom[3][37][35] = 2'b00;	 rom[3][38][35] = 2'b00;	 rom[3][39][35] = 2'b00;
 rom[3][0][36] = 2'b00;	 rom[3][1][36] = 2'b00;	 rom[3][2][36] = 2'b00;	 rom[3][3][36] = 2'b00;	 rom[3][4][36] = 2'b00;	 rom[3][5][36] = 2'b00;	 rom[3][6][36] = 2'b00;	 rom[3][7][36] = 2'b00;	 rom[3][8][36] = 2'b00;	 rom[3][9][36] = 2'b00;	 rom[3][10][36] = 2'b10;	 rom[3][11][36] = 2'b10;	 rom[3][12][36] = 2'b01;	 rom[3][13][36] = 2'b01;	 rom[3][14][36] = 2'b01;	 rom[3][15][36] = 2'b01;	 rom[3][16][36] = 2'b01;	 rom[3][17][36] = 2'b01;	 rom[3][18][36] = 2'b01;	 rom[3][19][36] = 2'b01;	 rom[3][20][36] = 2'b01;	 rom[3][21][36] = 2'b01;	 rom[3][22][36] = 2'b01;	 rom[3][23][36] = 2'b01;	 rom[3][24][36] = 2'b01;	 rom[3][25][36] = 2'b10;	 rom[3][26][36] = 2'b10;	 rom[3][27][36] = 2'b10;	 rom[3][28][36] = 2'b10;	 rom[3][29][36] = 2'b00;	 rom[3][30][36] = 2'b00;	 rom[3][31][36] = 2'b00;	 rom[3][32][36] = 2'b00;	 rom[3][33][36] = 2'b00;	 rom[3][34][36] = 2'b00;	 rom[3][35][36] = 2'b00;	 rom[3][36][36] = 2'b00;	 rom[3][37][36] = 2'b00;	 rom[3][38][36] = 2'b00;	 rom[3][39][36] = 2'b00;
 rom[3][0][37] = 2'b00;	 rom[3][1][37] = 2'b00;	 rom[3][2][37] = 2'b00;	 rom[3][3][37] = 2'b00;	 rom[3][4][37] = 2'b00;	 rom[3][5][37] = 2'b00;	 rom[3][6][37] = 2'b00;	 rom[3][7][37] = 2'b00;	 rom[3][8][37] = 2'b00;	 rom[3][9][37] = 2'b00;	 rom[3][10][37] = 2'b00;	 rom[3][11][37] = 2'b10;	 rom[3][12][37] = 2'b10;	 rom[3][13][37] = 2'b10;	 rom[3][14][37] = 2'b10;	 rom[3][15][37] = 2'b10;	 rom[3][16][37] = 2'b10;	 rom[3][17][37] = 2'b10;	 rom[3][18][37] = 2'b10;	 rom[3][19][37] = 2'b10;	 rom[3][20][37] = 2'b10;	 rom[3][21][37] = 2'b10;	 rom[3][22][37] = 2'b10;	 rom[3][23][37] = 2'b10;	 rom[3][24][37] = 2'b10;	 rom[3][25][37] = 2'b10;	 rom[3][26][37] = 2'b11;	 rom[3][27][37] = 2'b11;	 rom[3][28][37] = 2'b10;	 rom[3][29][37] = 2'b00;	 rom[3][30][37] = 2'b00;	 rom[3][31][37] = 2'b00;	 rom[3][32][37] = 2'b00;	 rom[3][33][37] = 2'b00;	 rom[3][34][37] = 2'b00;	 rom[3][35][37] = 2'b00;	 rom[3][36][37] = 2'b00;	 rom[3][37][37] = 2'b00;	 rom[3][38][37] = 2'b00;	 rom[3][39][37] = 2'b00;
 rom[3][0][38] = 2'b00;	 rom[3][1][38] = 2'b00;	 rom[3][2][38] = 2'b00;	 rom[3][3][38] = 2'b00;	 rom[3][4][38] = 2'b00;	 rom[3][5][38] = 2'b00;	 rom[3][6][38] = 2'b00;	 rom[3][7][38] = 2'b00;	 rom[3][8][38] = 2'b00;	 rom[3][9][38] = 2'b00;	 rom[3][10][38] = 2'b00;	 rom[3][11][38] = 2'b00;	 rom[3][12][38] = 2'b00;	 rom[3][13][38] = 2'b00;	 rom[3][14][38] = 2'b00;	 rom[3][15][38] = 2'b00;	 rom[3][16][38] = 2'b00;	 rom[3][17][38] = 2'b00;	 rom[3][18][38] = 2'b00;	 rom[3][19][38] = 2'b00;	 rom[3][20][38] = 2'b00;	 rom[3][21][38] = 2'b00;	 rom[3][22][38] = 2'b00;	 rom[3][23][38] = 2'b00;	 rom[3][24][38] = 2'b10;	 rom[3][25][38] = 2'b11;	 rom[3][26][38] = 2'b11;	 rom[3][27][38] = 2'b11;	 rom[3][28][38] = 2'b10;	 rom[3][29][38] = 2'b00;	 rom[3][30][38] = 2'b00;	 rom[3][31][38] = 2'b00;	 rom[3][32][38] = 2'b00;	 rom[3][33][38] = 2'b00;	 rom[3][34][38] = 2'b00;	 rom[3][35][38] = 2'b00;	 rom[3][36][38] = 2'b00;	 rom[3][37][38] = 2'b00;	 rom[3][38][38] = 2'b00;	 rom[3][39][38] = 2'b00;
 rom[3][0][39] = 2'b00;	 rom[3][1][39] = 2'b00;	 rom[3][2][39] = 2'b00;	 rom[3][3][39] = 2'b00;	 rom[3][4][39] = 2'b00;	 rom[3][5][39] = 2'b00;	 rom[3][6][39] = 2'b00;	 rom[3][7][39] = 2'b00;	 rom[3][8][39] = 2'b00;	 rom[3][9][39] = 2'b00;	 rom[3][10][39] = 2'b00;	 rom[3][11][39] = 2'b00;	 rom[3][12][39] = 2'b00;	 rom[3][13][39] = 2'b00;	 rom[3][14][39] = 2'b00;	 rom[3][15][39] = 2'b00;	 rom[3][16][39] = 2'b00;	 rom[3][17][39] = 2'b00;	 rom[3][18][39] = 2'b00;	 rom[3][19][39] = 2'b00;	 rom[3][20][39] = 2'b00;	 rom[3][21][39] = 2'b00;	 rom[3][22][39] = 2'b00;	 rom[3][23][39] = 2'b00;	 rom[3][24][39] = 2'b10;	 rom[3][25][39] = 2'b10;	 rom[3][26][39] = 2'b10;	 rom[3][27][39] = 2'b10;	 rom[3][28][39] = 2'b10;	 rom[3][29][39] = 2'b00;	 rom[3][30][39] = 2'b00;	 rom[3][31][39] = 2'b00;	 rom[3][32][39] = 2'b00;	 rom[3][33][39] = 2'b00;	 rom[3][34][39] = 2'b00;	 rom[3][35][39] = 2'b00;	 rom[3][36][39] = 2'b00;	 rom[3][37][39] = 2'b00;	 rom[3][38][39] = 2'b00;	 rom[3][39][39] = 2'b00;


end

assign data = en ? rom[dir][x][y] : 2'b00;

endmodule















